version https://git-lfs.github.com/spec/v1
oid sha256:caa2882567f6a82128169c0a5a9aaf8f109bcfab8277685b1de2f619d4dcb36c
size 11961

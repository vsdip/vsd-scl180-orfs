*  -------------------------------------- *
*  Filename: scl18fs120_supply_pins.cdl
*  Total subcircuits:  540
*  -------------------------------------- *
* Defining the default unit for both length and area
*.SCALE meter
*  -------------------------------------- *

.SUBCKT ad01d0 CO S  A B CI VDD VSS
MM28 VDD CI 7 VDD P l=0.191475u w=1.83u 
MM17 VDD A 7 VDD P l=0.18u w=1.37u 
MM27 13 CI 4 VDD P l=0.186301u w=1.314u 
MM26 13 B VDD VDD P l=0.18u w=1.26u 
MM25 VDD B 7 VDD P l=0.18u w=1.14u 
MM22 6 4 7 VDD P l=0.188502u w=1.235u 
MM20 6 CI 18 VDD P l=0.18u w=1.44u 
MM23 VDD B 17 VDD P l=0.18u w=1.44u 
MM21 17 A 18 VDD P l=0.18u w=1.44u 
MM19 19 A 4 VDD P l=0.18u w=1.24u 
MM24 VDD B 19 VDD P l=0.18u w=1.24u 
MM18 13 A VDD VDD P l=0.185865u w=1.33u 
MM16 VDD 4 CO VDD P l=0.18u w=0.85u 
MM15 S 6 VDD VDD P l=0.18u w=0.85u 
MM13 12 CI 4 VSS N l=0.186935u w=1.194u 
MM9 VSS B 12 VSS N l=0.18u w=1.23u 
MM14 9 CI VSS VSS N l=0.187312u w=1.198u 
MM8 6 4 9 VSS N l=0.185738u w=1.192u 
MM6 6 CI 15 VSS N l=0.18u w=1.12u 
MM12 VSS B 14 VSS N l=0.186935u w=1.194u 
MM7 14 A 15 VSS N l=0.18u w=1.12u 
MM5 4 A 16 VSS N l=0.18u w=1.12u 
MM10 VSS B 16 VSS N l=0.18u w=1.12u 
MM4 VSS A 12 VSS N l=0.186u w=1.3u 
MM11 9 B VSS VSS N l=0.186935u w=1.194u 
MM3 9 A VSS VSS N l=0.18u w=1.12u 
MM2 VSS 4 CO VSS N l=0.18u w=0.57u 
MM1 S 6 VSS VSS N l=0.18u w=0.57u 
.ENDS ad01d0

.SUBCKT ad01d1 CO S  A B CI VDD VSS
MM28 VDD CI 7 VDD P l=0.191475u w=1.83u 
MM17 VDD A 7 VDD P l=0.18u w=1.37u 
MM27 13 CI 4 VDD P l=0.186301u w=1.314u 
MM26 13 B VDD VDD P l=0.18u w=1.26u 
MM25 VDD B 7 VDD P l=0.18u w=1.14u 
MM22 6 4 7 VDD P l=0.188502u w=1.235u 
MM20 6 CI 18 VDD P l=0.18u w=1.44u 
MM23 VDD B 17 VDD P l=0.18u w=1.44u 
MM21 17 A 18 VDD P l=0.18u w=1.44u 
MM19 19 A 4 VDD P l=0.18u w=1.24u 
MM24 VDD B 19 VDD P l=0.18u w=1.24u 
MM18 13 A VDD VDD P l=0.185865u w=1.33u 
MM16 VDD 4 CO VDD P l=0.185099u w=1.624u 
MM15 VDD 6 S VDD P l=0.18u w=1.55u 
MM13 12 CI 4 VSS N l=0.186935u w=1.194u 
MM9 VSS B 12 VSS N l=0.18u w=1.23u 
MM14 9 CI VSS VSS N l=0.187312u w=1.198u 
MM8 6 4 9 VSS N l=0.185738u w=1.192u 
MM6 6 CI 15 VSS N l=0.18u w=1.12u 
MM12 VSS B 14 VSS N l=0.186935u w=1.194u 
MM7 14 A 15 VSS N l=0.18u w=1.12u 
MM5 4 A 16 VSS N l=0.18u w=1.12u 
MM10 VSS B 16 VSS N l=0.18u w=1.12u 
MM4 VSS A 12 VSS N l=0.186u w=1.3u 
MM11 9 B VSS VSS N l=0.186935u w=1.194u 
MM3 9 A VSS VSS N l=0.18u w=1.12u 
MM2 CO 4 VSS VSS N l=0.187569u w=1.094u 
MM1 VSS 6 S VSS N l=0.18u w=1.02u 
.ENDS ad01d1

.SUBCKT ad01d2 CO S  A B CI VDD VSS
MM32 13 B VDD VDD P l=0.18u w=1.26u 
MM17 13 CI 3 VDD P l=0.186301u w=1.314u 
MM29 VDD B 17 VDD P l=0.18u w=1.24u 
MM21 17 A 3 VDD P l=0.18u w=1.24u 
MM20 13 A VDD VDD P l=0.185865u w=1.33u 
MM30 VDD B 7 VDD P l=0.18u w=1.14u 
MM28 7 3 6 VDD P l=0.189575u w=1.247u 
MM19 VDD A 7 VDD P l=0.18u w=1.37u 
MM18 VDD CI 7 VDD P l=0.190759u w=1.818u 
MM31 VDD B 18 VDD P l=0.18u w=1.44u 
MM27 18 A 19 VDD P l=0.18u w=1.44u 
MM26 19 CI 6 VDD P l=0.18u w=1.44u 
MM23 VDD 6 S VDD P l=0.184436u w=1.542u 
MM22 VDD 6 S VDD P l=0.185328u w=1.554u 
MM25 VDD 3 CO VDD P l=0.185032u w=1.55u 
MM24 VDD 3 CO VDD P l=0.18u w=1.48u 
MM13 VSS B 12 VSS N l=0.18u w=1.2u 
MM1 12 CI 3 VSS N l=0.187113u w=1.164u 
MM14 VSS B 14 VSS N l=0.18u w=1.09u 
MM5 3 A 14 VSS N l=0.18u w=1.09u 
MM4 VSS A 12 VSS N l=0.186499u w=1.274u 
MM15 9 B VSS VSS N l=0.187113u w=1.164u 
MM3 9 A VSS VSS N l=0.18u w=1.09u 
MM12 6 3 9 VSS N l=0.185937u w=1.152u 
MM2 9 CI VSS VSS N l=0.187113u w=1.164u 
MM16 VSS B 15 VSS N l=0.189652u w=1.237u 
MM11 15 A 16 VSS N l=0.18u w=1.09u 
MM10 6 CI 16 VSS N l=0.18u w=1.09u 
MM7 VSS 6 S VSS N l=0.186998u w=1.046u 
MM6 VSS 6 S VSS N l=0.18u w=0.98u 
MM9 VSS 3 CO VSS N l=0.186693u w=1.022u 
MM8 VSS 3 CO VSS N l=0.18u w=0.96u 
.ENDS ad01d2

.SUBCKT adiode   I VDD VSS
D1      VSS   I DN  462.4000F 2.7200U
D2      I   VDD DP  462.4000F 2.7200U
.ENDS adiode

.SUBCKT adp1d0 CO P S  A B CI VDD VSS
MM38 24 2 6 VDD P l=0.18u w=1.54u 
MM36 6 A 23 VDD P l=0.18427u w=1.602u 
MM37 VDD B 23 VDD P l=0.18513u w=1.614u 
MM35 24 5 VDD VDD P l=0.18u w=1.54u 
MM34 P 6 VDD VDD P l=0.18u w=1.54u 
MM29 CO 9 VDD VDD P l=0.18u w=0.56u 
MM33 14 B VDD VDD P l=0.186301u w=1.314u 
MM31 9 7 14 VDD P l=0.18u w=1.24u 
MM30 9 CI 14 VDD P l=0.186301u w=1.314u 
MM32 VDD A 14 VDD P l=0.18u w=1.24u 
MM28 VDD B 5 VDD P l=0.18u w=0.55u 
MM27 VDD A 2 VDD P l=0.18u w=0.55u 
MM25 25 7 11 VDD P l=0.18u w=1.54u 
MM22 11 6 26 VDD P l=0.185398u w=1.534u 
MM24 S 11 VDD VDD P l=0.184845u w=1.61u 
MM23 25 CI VDD VDD P l=0.18u w=1.54u 
MM26 VDD 10 26 VDD P l=0.185398u w=1.534u 
MM21 VDD 6 7 VDD P l=0.18u w=0.58u 
MM20 10 CI VDD VDD P l=0.18u w=0.63u 
MM19 17 2 6 VSS N l=0.18u w=0.81u 
MM18 VSS B 17 VSS N l=0.18u w=0.81u 
MM17 5 B VSS VSS N l=0.18u w=0.48u 
MM16 18 A VSS VSS N l=0.18u w=0.81u 
MM15 18 5 6 VSS N l=0.18u w=0.81u 
MM14 VSS 6 P VSS N l=0.18u w=1.54u 
MM12 2 A VSS VSS N l=0.18u w=0.42u 
MM13 19 B VSS VSS N l=0.18u w=0.88u 
MM11 9 A 19 VSS N l=0.18u w=0.88u 
MM10 20 7 9 VSS N l=0.18u w=0.88u 
MM9 20 CI VSS VSS N l=0.18u w=0.88u 
MM8 CO 9 VSS VSS N l=0.18u w=0.46u 
MM7 10 CI VSS VSS N l=0.18u w=0.48u 
MM6 21 10 VSS VSS N l=0.18u w=0.74u 
MM5 21 7 11 VSS N l=0.18u w=0.74u 
MM4 S 11 VSS VSS N l=0.187222u w=1.08u 
MM2 7 6 VSS VSS N l=0.18u w=0.5u 
MM1 11 6 22 VSS N l=0.18u w=0.74u 
MM3 22 CI VSS VSS N l=0.18u w=0.74u 
.ENDS adp1d0

.SUBCKT adp1d1 CO P S  A B CI VDD VSS
MM38 24 2 6 VDD P l=0.18u w=1.54u 
MM36 6 A 23 VDD P l=0.18427u w=1.602u 
MM37 VDD B 23 VDD P l=0.18513u w=1.614u 
MM35 24 5 VDD VDD P l=0.18u w=1.54u 
MM34 P 6 VDD VDD P l=0.18u w=1.54u 
MM33 14 B VDD VDD P l=0.186254u w=1.324u 
MM31 9 7 14 VDD P l=0.18u w=1.17u 
MM32 VDD A 14 VDD P l=0.18u w=1.17u 
MM30 9 CI 14 VDD P l=0.186656u w=1.244u 
MM29 CO 9 VDD VDD P l=0.185562u w=1.316u 
MM28 VDD B 5 VDD P l=0.18u w=0.55u 
MM27 VDD A 2 VDD P l=0.18u w=0.55u 
MM25 25 7 11 VDD P l=0.18u w=1.54u 
MM22 11 6 26 VDD P l=0.185398u w=1.534u 
MM24 S 11 VDD VDD P l=0.184845u w=1.61u 
MM23 25 CI VDD VDD P l=0.18u w=1.54u 
MM26 VDD 10 26 VDD P l=0.185398u w=1.534u 
MM21 VDD 6 7 VDD P l=0.18u w=0.58u 
MM20 10 CI VDD VDD P l=0.18u w=0.65u 
MM19 17 2 6 VSS N l=0.18u w=0.81u 
MM18 VSS B 17 VSS N l=0.18u w=0.81u 
MM17 5 B VSS VSS N l=0.18u w=0.48u 
MM16 18 A VSS VSS N l=0.18u w=0.81u 
MM15 18 5 6 VSS N l=0.18u w=0.81u 
MM14 VSS 6 P VSS N l=0.18u w=1.54u 
MM12 2 A VSS VSS N l=0.18u w=0.42u 
MM13 19 B VSS VSS N l=0.18u w=0.88u 
MM11 9 A 19 VSS N l=0.18u w=0.88u 
MM10 20 7 9 VSS N l=0.18u w=0.88u 
MM9 20 CI VSS VSS N l=0.18u w=0.88u 
MM8 CO 9 VSS VSS N l=0.185978u w=1.626u 
MM7 10 CI VSS VSS N l=0.18u w=0.48u 
MM6 21 10 VSS VSS N l=0.18u w=0.74u 
MM5 21 7 11 VSS N l=0.18u w=0.74u 
MM4 S 11 VSS VSS N l=0.187222u w=1.08u 
MM2 7 6 VSS VSS N l=0.18u w=0.5u 
MM1 11 6 22 VSS N l=0.18u w=0.74u 
MM3 22 CI VSS VSS N l=0.18u w=0.74u 
.ENDS adp1d1

.SUBCKT adp1d2 CO P S  A B CI VDD VSS
MM40 24 2 6 VDD P l=0.18u w=1.54u 
MM38 6 A 23 VDD P l=0.18427u w=1.602u 
MM39 VDD B 23 VDD P l=0.18513u w=1.614u 
MM37 24 5 VDD VDD P l=0.18u w=1.54u 
MM36 P 6 VDD VDD P l=0.18u w=1.54u 
MM35 VDD B 5 VDD P l=0.18u w=0.55u 
MM34 VDD A 2 VDD P l=0.18u w=0.55u 
MM33 14 B VDD VDD P l=0.186254u w=1.324u 
MM31 9 7 14 VDD P l=0.18u w=1.17u 
MM32 VDD A 14 VDD P l=0.18u w=1.17u 
MM30 9 CI 14 VDD P l=0.186656u w=1.244u 
MM29 CO 9 VDD VDD P l=0.186449u w=1.284u 
MM28 CO 9 VDD VDD P l=0.18u w=1.21u 
MM26 25 7 11 VDD P l=0.18u w=1.54u 
MM23 11 6 26 VDD P l=0.185398u w=1.534u 
MM25 S 11 VDD VDD P l=0.184845u w=1.61u 
MM24 25 CI VDD VDD P l=0.18u w=1.54u 
MM27 VDD 10 26 VDD P l=0.185398u w=1.534u 
MM22 VDD 6 7 VDD P l=0.18u w=0.58u 
MM21 10 CI VDD VDD P l=0.18u w=0.65u 
MM20 17 2 6 VSS N l=0.18u w=0.81u 
MM19 VSS B 17 VSS N l=0.18u w=0.81u 
MM18 5 B VSS VSS N l=0.18u w=0.48u 
MM17 18 A VSS VSS N l=0.18u w=0.81u 
MM16 6 5 18 VSS N l=0.18u w=0.81u 
MM15 VSS 6 P VSS N l=0.18u w=1.54u 
MM13 2 A VSS VSS N l=0.18u w=0.45u 
MM14 19 B VSS VSS N l=0.18u w=0.91u 
MM12 9 A 19 VSS N l=0.18u w=0.91u 
MM11 20 7 9 VSS N l=0.18u w=0.91u 
MM10 20 CI VSS VSS N l=0.18u w=0.91u 
MM9 CO 9 VSS VSS N l=0.188196u w=1.186u 
MM8 CO 9 VSS VSS N l=0.18u w=1.1u 
MM7 10 CI VSS VSS N l=0.18u w=0.48u 
MM6 21 10 VSS VSS N l=0.18u w=0.74u 
MM5 21 7 11 VSS N l=0.18u w=0.74u 
MM4 S 11 VSS VSS N l=0.187222u w=1.08u 
MM2 7 6 VSS VSS N l=0.18u w=0.5u 
MM1 22 6 11 VSS N l=0.18u w=0.74u 
MM3 22 CI VSS VSS N l=0.18u w=0.74u 
.ENDS adp1d2

.SUBCKT ah01d0 CO S  A B VDD VSS
MM14 VDD 2 5 VDD P l=0.18u w=0.57u 
MM13 5 A 11 VDD P l=0.18u w=1.14u 
MM12 VDD B 11 VDD P l=0.18u w=1.14u 
MM11 VDD 2 CO VDD P l=0.18u w=0.72u 
MM10 VDD 5 S VDD P l=0.18u w=0.72u 
MM9 VDD A 2 VDD P l=0.18u w=0.57u 
MM8 VDD B 2 VDD P l=0.18u w=0.57u 
MM7 2 A 10 VSS N l=0.18u w=0.82u 
MM6 9 A VSS VSS N l=0.18u w=0.57u 
MM5 5 2 9 VSS N l=0.18u w=0.72u 
MM3 9 B VSS VSS N l=0.18u w=0.82u 
MM4 VSS B 10 VSS N l=0.18u w=0.82u 
MM2 CO 2 VSS VSS N l=0.18u w=0.5u 
MM1 S 5 VSS VSS N l=0.18u w=0.5u 
.ENDS ah01d0

.SUBCKT ah01d1 CO S  A B VDD VSS
MM14 VDD 2 5 VDD P l=0.18u w=0.57u 
MM13 5 A 11 VDD P l=0.18u w=1.14u 
MM12 VDD B 11 VDD P l=0.18u w=1.14u 
MM11 CO 2 VDD VDD P l=0.184584u w=1.492u 
MM10 S 5 VDD VDD P l=0.1852u w=1.5u 
MM9 VDD A 2 VDD P l=0.18u w=0.57u 
MM8 VDD B 2 VDD P l=0.18u w=0.57u 
MM7 5 2 9 VSS N l=0.18u w=0.72u 
MM5 9 A VSS VSS N l=0.18u w=0.57u 
MM3 VSS B 9 VSS N l=0.18u w=0.82u 
MM6 2 A 10 VSS N l=0.18u w=0.82u 
MM4 VSS B 10 VSS N l=0.18u w=0.82u 
MM2 CO 2 VSS VSS N l=0.18u w=0.95u 
MM1 S 5 VSS VSS N l=0.18u w=0.95u 
.ENDS ah01d1

.SUBCKT ah01d2 CO S  A B VDD VSS
MM18 VDD 2 5 VDD P l=0.18u w=0.57u 
MM17 11 A 5 VDD P l=0.18u w=1.14u 
MM16 VDD B 11 VDD P l=0.18u w=1.14u 
MM15 CO 2 VDD VDD P l=0.185505u w=1.504u 
MM14 CO 2 VDD VDD P l=0.18u w=1.43u 
MM13 VDD 5 S VDD P l=0.1852u w=1.5u 
MM12 S 5 VDD VDD P l=0.18u w=1.43u 
MM11 VDD A 2 VDD P l=0.18u w=0.57u 
MM10 VDD B 2 VDD P l=0.18u w=0.57u 
MM9 9 2 5 VSS N l=0.18u w=0.72u 
MM7 9 A VSS VSS N l=0.18u w=0.57u 
MM5 9 B VSS VSS N l=0.18u w=0.82u 
MM8 2 A 10 VSS N l=0.18u w=0.82u 
MM6 VSS B 10 VSS N l=0.18u w=0.82u 
MM4 VSS 2 CO VSS N l=0.18u w=0.95u 
MM3 VSS 2 CO VSS N l=0.18u w=0.95u 
MM2 VSS 5 S VSS N l=0.18u w=0.95u 
MM1 VSS 5 S VSS N l=0.18u w=0.95u 
.ENDS ah01d2

.SUBCKT an02d0 Z  A1 A2 VDD VSS
MM5 VDD 3 Z VDD P l=0.18u w=0.74u 
MM6 VDD A2 3 VDD P l=0.18u w=0.88u 
MM4 VDD A1 3 VDD P l=0.18u w=0.88u 
MM2 VSS 3 Z VSS N l=0.18u w=0.5u 
MM3 7 A2 VSS VSS N l=0.18u w=0.88u 
MM1 7 A1 3 VSS N l=0.18u w=0.88u 
.ENDS an02d0

.SUBCKT an02d1 Z  A1 A2 VDD VSS
MM5 VDD 3 Z VDD P l=0.18u w=1.48u 
MM6 VDD A2 3 VDD P l=0.18u w=0.88u 
MM4 VDD A1 3 VDD P l=0.18u w=0.88u 
MM2 Z 3 VSS VSS N l=0.18u w=1u 
MM3 7 A2 VSS VSS N l=0.18u w=0.88u 
MM1 7 A1 3 VSS N l=0.18u w=0.88u 
.ENDS an02d1

.SUBCKT an02d2 Z  A1 A2 VDD VSS
MM8 VDD 2 Z VDD P l=0.184937u w=1.58u 
MM7 VDD 2 Z VDD P l=0.18u w=1.51u 
MM6 VDD A2 2 VDD P l=0.18u w=0.7u 
MM5 VDD A1 2 VDD P l=0.18u w=0.7u 
MM4 Z 2 VSS VSS N l=0.187864u w=1.236u 
MM3 Z 2 VSS VSS N l=0.18u w=1.15u 
MM2 VSS A2 7 VSS N l=0.18u w=0.7u 
MM1 7 A1 2 VSS N l=0.18u w=0.7u 
.ENDS an02d2

.SUBCKT an02d4 Z  A1 A2 VDD VSS
MM10 VDD 2 Z VDD P l=0.184012u w=2.064u 
MM9 VDD 2 Z VDD P l=0.18u w=1.99u 
MM8 VDD 2 Z VDD P l=0.184012u w=2.064u 
MM7 2 A2 VDD VDD P l=0.18u w=1.4u 
MM6 2 A1 VDD VDD P l=0.184993u w=1.466u 
MM5 VSS 2 Z VSS N l=0.186454u w=1.506u 
MM4 VSS 2 Z VSS N l=0.186152u w=1.502u 
MM3 VSS 2 Z VSS N l=0.18u w=1.42u 
MM2 VSS A2 7 VSS N l=0.18u w=0.7u 
MM1 7 A1 2 VSS N l=0.18u w=0.7u 
.ENDS an02d4

.SUBCKT an03d0 Z  A1 A2 A3 VDD VSS
MM7 VDD 3 Z VDD P l=0.18u w=0.7u 
MM8 3 A3 VDD VDD P l=0.18u w=0.78u 
MM6 3 A2 VDD VDD P l=0.18u w=0.78u 
MM5 3 A1 VDD VDD P l=0.18u w=0.78u 
MM3 VSS 3 Z VSS N l=0.18u w=0.62u 
MM4 VSS A3 8 VSS N l=0.18u w=0.8u 
MM2 8 A2 9 VSS N l=0.18u w=0.8u 
MM1 3 A1 9 VSS N l=0.18u w=0.8u 
.ENDS an03d0

.SUBCKT an03d1 Z  A1 A2 A3 VDD VSS
MM7 VDD 3 Z VDD P l=0.185417u w=1.44u 
MM8 3 A3 VDD VDD P l=0.18u w=0.78u 
MM6 3 A2 VDD VDD P l=0.18u w=0.78u 
MM5 3 A1 VDD VDD P l=0.18u w=0.78u 
MM3 VSS 3 Z VSS N l=0.18542u w=1.262u 
MM4 VSS A3 8 VSS N l=0.18u w=0.8u 
MM2 8 A2 9 VSS N l=0.18u w=0.8u 
MM1 3 A1 9 VSS N l=0.18u w=0.8u 
.ENDS an03d1

.SUBCKT an03d2 Z  A1 A2 A3 VDD VSS
MM7 3 A1 VDD VDD P l=0.18u w=0.78u 
MM9 VDD 3 Z VDD P l=0.185417u w=1.44u 
MM8 Z 3 VDD VDD P l=0.18u w=1.37u 
MM10 3 A3 VDD VDD P l=0.18u w=0.78u 
MM6 3 A2 VDD VDD P l=0.18u w=0.78u 
MM4 VSS 3 Z VSS N l=0.186142u w=1.27u 
MM3 VSS 3 Z VSS N l=0.18u w=1.2u 
MM2 3 A1 9 VSS N l=0.18u w=0.8u 
MM5 VSS A3 8 VSS N l=0.18u w=0.8u 
MM1 8 A2 9 VSS N l=0.18u w=0.8u 
.ENDS an03d2

.SUBCKT an03d4 Z  A1 A2 A3 VDD VSS
MM12 VDD 2 Z VDD P l=0.183786u w=2.06u 
MM11 Z 2 VDD VDD P l=0.18u w=1.99u 
MM10 Z 2 VDD VDD P l=0.183786u w=2.06u 
MM9 VDD A3 2 VDD P l=0.18u w=1.51u 
MM8 VDD A2 2 VDD P l=0.18u w=1.51u 
MM7 VDD A1 2 VDD P l=0.18u w=1.51u 
MM6 VSS 2 Z VSS N l=0.185067u w=1.634u 
MM5 VSS 2 Z VSS N l=0.18u w=1.56u 
MM4 VSS 2 Z VSS N l=0.18u w=1.56u 
MM3 8 A3 VSS VSS N l=0.18u w=1.16u 
MM2 9 A2 8 VSS N l=0.18u w=1.16u 
MM1 9 A1 2 VSS N l=0.18u w=1.16u 
.ENDS an03d4

.SUBCKT an04d0 Z  A1 A2 A3 A4 VDD VSS
MM10 VDD 2 Z VDD P l=0.18u w=0.63u 
MM9 VDD A4 2 VDD P l=0.18u w=0.87u 
MM8 VDD A3 2 VDD P l=0.18u w=0.87u 
MM7 VDD A2 2 VDD P l=0.18u w=0.87u 
MM6 VDD A1 2 VDD P l=0.18u w=0.87u 
MM5 VSS 2 Z VSS N l=0.18u w=0.5u 
MM4 9 A4 VSS VSS N l=0.18u w=0.9u 
MM3 9 A3 10 VSS N l=0.18u w=0.9u 
MM2 11 A2 10 VSS N l=0.18u w=0.9u 
MM1 2 A1 11 VSS N l=0.18u w=0.9u 
.ENDS an04d0

.SUBCKT an04d1 Z  A1 A2 A3 A4 VDD VSS
MM9 Z 3 VDD VDD P l=0.18u w=1.26u 
MM10 VDD A4 3 VDD P l=0.18u w=0.87u 
MM8 VDD A3 3 VDD P l=0.18u w=0.87u 
MM7 VDD A2 3 VDD P l=0.18u w=0.87u 
MM6 VDD A1 3 VDD P l=0.18u w=0.87u 
MM4 Z 3 VSS VSS N l=0.18u w=1u 
MM5 VSS A4 9 VSS N l=0.18u w=0.9u 
MM3 10 A3 9 VSS N l=0.18u w=0.9u 
MM2 10 A2 11 VSS N l=0.18u w=0.9u 
MM1 3 A1 11 VSS N l=0.18u w=0.9u 
.ENDS an04d1

.SUBCKT an04d2 Z  A1 A2 A3 A4 VDD VSS
MM11 Z 3 VDD VDD P l=0.18u w=1.26u 
MM10 Z 3 VDD VDD P l=0.18u w=1.26u 
MM12 VDD A4 3 VDD P l=0.18u w=0.87u 
MM9 VDD A3 3 VDD P l=0.18u w=0.87u 
MM8 VDD A2 3 VDD P l=0.18u w=0.87u 
MM7 VDD A1 3 VDD P l=0.18u w=0.87u 
MM5 Z 3 VSS VSS N l=0.18u w=1u 
MM4 VSS 3 Z VSS N l=0.18u w=1u 
MM6 VSS A4 9 VSS N l=0.18u w=0.9u 
MM3 10 A3 9 VSS N l=0.18u w=0.9u 
MM2 10 A2 11 VSS N l=0.18u w=0.9u 
MM1 3 A1 11 VSS N l=0.18u w=0.9u 
.ENDS an04d2

.SUBCKT an04d4 Z  A1 A2 A3 A4 VDD VSS
MM13 Z 3 VDD VDD P l=0.184457u w=1.75u 
MM12 VDD 3 Z VDD P l=0.184721u w=1.754u 
MM11 VDD 3 Z VDD P l=0.18u w=1.68u 
MM14 VDD A4 3 VDD P l=0.18u w=1.4u 
MM10 3 A3 VDD VDD P l=0.18u w=1.4u 
MM9 3 A2 VDD VDD P l=0.18u w=1.4u 
MM8 3 A1 VDD VDD P l=0.18u w=1.4u 
MM6 Z 3 VSS VSS N l=0.185856u w=1.414u 
MM5 Z 3 VSS VSS N l=0.18u w=1.34u 
MM4 Z 3 VSS VSS N l=0.18u w=1.34u 
MM7 VSS A4 9 VSS N l=0.18u w=1.17u 
MM3 10 A3 9 VSS N l=0.18u w=1.17u 
MM2 11 A2 10 VSS N l=0.18u w=1.17u 
MM1 11 A1 3 VSS N l=0.18u w=1.17u 
.ENDS an04d4

.SUBCKT an12d1 Z  A1 A2 VDD VSS
MM7 Z 3 VDD VDD P l=0.184937u w=1.58u 
MM6 5 A1 VDD VDD P l=0.18u w=0.62u 
MM8 VDD A2 3 VDD P l=0.18u w=0.87u 
MM5 VDD 5 3 VDD P l=0.18u w=0.87u 
MM3 Z 3 VSS VSS N l=0.185738u w=1.192u 
MM4 8 A2 VSS VSS N l=0.18u w=0.9u 
MM2 8 5 3 VSS N l=0.18u w=0.9u 
MM1 5 A1 VSS VSS N l=0.18u w=0.48u 
.ENDS an12d1

.SUBCKT an12d2 Z  A1 A2 VDD VSS
MM9 VDD 3 Z VDD P l=0.184937u w=1.58u 
MM8 Z 3 VDD VDD P l=0.18u w=1.51u 
MM7 5 A1 VDD VDD P l=0.18u w=0.62u 
MM10 VDD A2 3 VDD P l=0.18u w=0.87u 
MM6 VDD 5 3 VDD P l=0.18u w=0.87u 
MM4 VSS 3 Z VSS N l=0.185738u w=1.192u 
MM3 VSS 3 Z VSS N l=0.18u w=1.13u 
MM5 8 A2 VSS VSS N l=0.18u w=0.9u 
MM2 8 5 3 VSS N l=0.18u w=0.9u 
MM1 5 A1 VSS VSS N l=0.18u w=0.48u 
.ENDS an12d2

.SUBCKT an12d4 Z  A1 A2 VDD VSS
MM12 Z 2 VDD VDD P l=0.183786u w=2.06u 
MM11 Z 2 VDD VDD P l=0.18u w=1.99u 
MM10 Z 2 VDD VDD P l=0.183786u w=2.06u 
MM9 5 A1 VDD VDD P l=0.18u w=0.78u 
MM8 VDD A2 2 VDD P l=0.18u w=1.41u 
MM7 VDD 5 2 VDD P l=0.18u w=1.41u 
MM6 VSS 2 Z VSS N l=0.185342u w=1.46u 
MM5 VSS 2 Z VSS N l=0.184711u w=1.452u 
MM4 VSS 2 Z VSS N l=0.18u w=1.39u 
MM3 8 A2 VSS VSS N l=0.18u w=1.16u 
MM2 8 5 2 VSS N l=0.18u w=1.16u 
MM1 5 A1 VSS VSS N l=0.18u w=0.48u 
.ENDS an12d4

.SUBCKT aoi211d1 ZN  A B C1 C2 VDD VSS
MM8 10 B 7 VDD P l=0.184766u w=1.536u 
MM7 7 C1 VDD VDD P l=0.186096u w=1.122u 
MM6 7 C2 VDD VDD P l=0.186903u w=1.13u 
MM5 10 A ZN VDD P l=0.184766u w=1.536u 
MM4 VSS B ZN VSS N l=0.188163u w=1.132u 
MM3 9 C1 ZN VSS N l=0.18u w=1.05u 
MM2 VSS C2 9 VSS N l=0.188163u w=1.132u 
MM1 VSS A ZN VSS N l=0.18u w=0.99u 
.ENDS aoi211d1

.SUBCKT aoi211d2 ZN  A B C1 C2 VDD VSS
MM14 6 A 12 VDD P l=0.18u w=1.47u 
MM13 10 B 12 VDD P l=0.18u w=1.47u 
MM12 VDD C1 10 VDD P l=0.186096u w=1.122u 
MM11 10 C2 VDD VDD P l=0.186903u w=1.13u 
MM10 7 6 VDD VDD P l=0.185787u w=1.182u 
MM9 ZN 7 VDD VDD P l=0.184043u w=1.692u 
MM8 ZN 7 VDD VDD P l=0.18u w=1.63u 
MM7 6 A VSS VSS N l=0.18u w=0.99u 
MM6 6 B VSS VSS N l=0.188782u w=1.141u 
MM5 11 C1 6 VSS N l=0.18u w=1.05u 
MM4 11 C2 VSS VSS N l=0.188163u w=1.132u 
MM3 VSS 6 7 VSS N l=0.18u w=0.84u 
MM2 VSS 7 ZN VSS N l=0.188585u w=1.279u 
MM1 VSS 7 ZN VSS N l=0.18u w=1.18u 
.ENDS aoi211d2

.SUBCKT aoi211d4 ZN  A B C1 C2 VDD VSS
MM16 3 2 VDD VDD P l=0.18u w=1.66u 
MM15 VDD 3 ZN VDD P l=0.183786u w=2.06u 
MM14 ZN 3 VDD VDD P l=0.184012u w=2.064u 
MM13 ZN 3 VDD VDD P l=0.18u w=1.99u 
MM12 2 A 12 VDD P l=0.18u w=1.47u 
MM11 12 B 10 VDD P l=0.18u w=1.47u 
MM10 VDD C1 10 VDD P l=0.186096u w=1.122u 
MM9 10 C2 VDD VDD P l=0.186903u w=1.13u 
MM8 3 2 VSS VSS N l=0.18u w=1.16u 
MM6 VSS 3 ZN VSS N l=0.184643u w=1.68u 
MM7 ZN 3 VSS VSS N l=0.184917u w=1.684u 
MM5 ZN 3 VSS VSS N l=0.18u w=1.61u 
MM4 2 A VSS VSS N l=0.185922u w=1.236u 
MM3 2 B VSS VSS N l=0.18u w=1.05u 
MM2 11 C1 2 VSS N l=0.18u w=1.05u 
MM1 11 C2 VSS VSS N l=0.186964u w=1.12u 
.ENDS aoi211d4

.SUBCKT aoi21d1 ZN  A B1 B2 VDD VSS
MM5 5 B2 VDD VDD P l=0.18624u w=1.25u 
MM6 5 B1 VDD VDD P l=0.185507u w=1.242u 
MM4 ZN A 5 VDD P l=0.18u w=1.18u 
MM3 ZN B1 8 VSS N l=0.18u w=1.05u 
MM2 VSS B2 8 VSS N l=0.188163u w=1.132u 
MM1 ZN A VSS VSS N l=0.188556u w=1.136u 
.ENDS aoi21d1

.SUBCKT aoi21d2 ZN  A B1 B2 VDD VSS
MM12 3 2 VDD VDD P l=0.185507u w=1.242u 
MM11 ZN 3 VDD VDD P l=0.183838u w=1.782u 
MM10 VDD 3 ZN VDD P l=0.183838u w=1.782u 
MM9 2 A 9 VDD P l=0.18u w=1.18u 
MM8 VDD B1 9 VDD P l=0.185507u w=1.242u 
MM7 VDD B2 9 VDD P l=0.18624u w=1.25u 
MM6 VSS A 2 VSS N l=0.188632u w=1.126u 
MM5 2 B1 10 VSS N l=0.18u w=1.04u 
MM4 VSS B2 10 VSS N l=0.188632u w=1.126u 
MM3 VSS 2 3 VSS N l=0.18u w=0.88u 
MM2 VSS 3 ZN VSS N l=0.187386u w=1.316u 
MM1 ZN 3 VSS VSS N l=0.18u w=1.23u 
.ENDS aoi21d2

.SUBCKT aoi21d4 ZN  A B1 B2 VDD VSS
MM14 VDD 2 3 VDD P l=0.18u w=0.89u 
MM13 ZN 3 VDD VDD P l=0.183786u w=2.06u 
MM12 VDD 3 ZN VDD P l=0.184012u w=2.064u 
MM11 VDD 3 ZN VDD P l=0.18u w=1.99u 
MM10 9 B1 VDD VDD P l=0.18u w=1.14u 
MM8 9 A 2 VDD P l=0.18u w=0.82u 
MM9 9 B2 VDD VDD P l=0.186446u w=1.21u 
MM7 3 2 VSS VSS N l=0.18u w=0.42u 
MM5 ZN 3 VSS VSS N l=0.184643u w=1.68u 
MM6 ZN 3 VSS VSS N l=0.184917u w=1.684u 
MM4 ZN 3 VSS VSS N l=0.18u w=1.61u 
MM3 2 B1 10 VSS N l=0.18u w=1.17u 
MM1 2 A VSS VSS N l=0.18u w=0.43u 
MM2 VSS B2 10 VSS N l=0.18629u w=1.24u 
.ENDS aoi21d4

.SUBCKT aoi221d1 ZN  A B1 B2 C1 C2 VDD VSS
MM7 8 B1 9 VDD P l=0.18u w=1.38u 
MM10 VDD C2 8 VDD P l=0.184815u w=1.62u 
MM9 8 C1 VDD VDD P l=0.18u w=1.55u 
MM8 8 B2 9 VDD P l=0.185132u w=1.52u 
MM6 ZN A 9 VDD P l=0.186541u w=1.486u 
MM5 ZN C2 11 VSS N l=0.18u w=0.98u 
MM4 11 C1 VSS VSS N l=0.18u w=0.98u 
MM3 12 B2 VSS VSS N l=0.18u w=0.98u 
MM2 12 B1 ZN VSS N l=0.18u w=1u 
MM1 ZN A VSS VSS N l=0.18u w=1u 
.ENDS aoi221d1

.SUBCKT aoi221d2 ZN  A B1 B2 C1 C2 VDD VSS
MM16 9 C1 VDD VDD P l=0.184019u w=1.702u 
MM14 9 B2 12 VDD P l=0.18u w=1.55u 
MM15 VDD C2 9 VDD P l=0.184019u w=1.702u 
MM13 9 B1 12 VDD P l=0.184815u w=1.62u 
MM12 7 6 VDD VDD P l=0.184286u w=1.82u 
MM11 ZN 7 VDD VDD P l=0.184286u w=1.82u 
MM10 ZN 7 VDD VDD P l=0.18u w=1.75u 
MM9 12 A 6 VDD P l=0.186419u w=1.561u 
MM8 13 C1 6 VSS N l=0.18u w=0.98u 
MM7 7 6 VSS VSS N l=0.187952u w=1.66u 
MM6 VSS 7 ZN VSS N l=0.188221u w=1.664u 
MM5 ZN 7 VSS VSS N l=0.18u w=1.54u 
MM4 13 C2 VSS VSS N l=0.18u w=0.98u 
MM3 VSS A 6 VSS N l=0.189091u w=1.155u 
MM1 14 B1 6 VSS N l=0.18u w=1.06u 
MM2 VSS B2 14 VSS N l=0.18u w=1.06u 
.ENDS aoi221d2

.SUBCKT aoi221d4 ZN  A B1 B2 C1 C2 VDD VSS
MM20 VDD C2 9 VDD P l=0.18u w=1.64u 
MM19 VDD C1 9 VDD P l=0.184831u w=1.714u 
MM18 9 B2 12 VDD P l=0.18u w=1.55u 
MM17 9 B1 12 VDD P l=0.184815u w=1.62u 
MM16 7 6 VDD VDD P l=0.184286u w=1.82u 
MM14 ZN 7 VDD VDD P l=0.18u w=1.52u 
MM13 ZN 7 VDD VDD P l=0.185482u w=1.598u 
MM15 ZN 7 VDD VDD P l=0.184324u w=1.582u 
MM12 VDD 7 ZN VDD P l=0.18u w=1.75u 
MM11 12 A 6 VDD P l=0.185065u w=1.54u 
MM9 7 6 VSS VSS N l=0.188354u w=1.58u 
MM7 VSS 7 ZN VSS N l=0.184797u w=1.526u 
MM6 VSS 7 ZN VSS N l=0.18u w=1.46u 
MM8 VSS 7 ZN VSS N l=0.185098u w=1.53u 
MM5 ZN 7 VSS VSS N l=0.18u w=1.46u 
MM10 13 C2 VSS VSS N l=0.18u w=0.98u 
MM4 13 C1 6 VSS N l=0.18u w=0.98u 
MM3 VSS A 6 VSS N l=0.189091u w=1.155u 
MM1 14 B1 6 VSS N l=0.18u w=1.06u 
MM2 VSS B2 14 VSS N l=0.18u w=1.06u 
.ENDS aoi221d4

.SUBCKT aoi2222d1 ZN  A1 A2 B1 B2 C1 C2 D1 D2 VDD VSS
MM22 4 2 VDD VDD P l=0.18u w=1.09u 
MM21 VDD 3 4 VDD P l=0.185937u w=1.152u 
MM20 ZN 4 VDD VDD P l=0.184173u w=1.984u 
MM19 3 C2 14 VDD P l=0.185532u w=1.41u 
MM18 3 C1 14 VDD P l=0.18u w=1.34u 
MM17 VDD D1 14 VDD P l=0.184432u w=1.76u 
MM16 VDD D2 14 VDD P l=0.18u w=1.69u 
MM15 16 B2 VDD VDD P l=0.18u w=1.72u 
MM14 16 B1 VDD VDD P l=0.184358u w=1.79u 
MM13 16 A1 2 VDD P l=0.18u w=1.42u 
MM12 16 A2 2 VDD P l=0.185235u w=1.49u 
MM10 17 3 4 VSS N l=0.18u w=1.17u 
MM11 17 2 VSS VSS N l=0.18u w=1.17u 
MM9 ZN 4 VSS VSS N l=0.18u w=1.19u 
MM8 18 C2 VSS VSS N l=0.18u w=0.72u 
MM7 18 C1 3 VSS N l=0.18u w=0.72u 
MM6 3 D1 19 VSS N l=0.18u w=0.87u 
MM5 VSS D2 19 VSS N l=0.18u w=0.87u 
MM4 20 B2 VSS VSS N l=0.18u w=1u 
MM3 20 B1 2 VSS N l=0.186867u w=1.066u 
MM2 2 A1 21 VSS N l=0.18u w=0.72u 
MM1 VSS A2 21 VSS N l=0.18u w=0.72u 
.ENDS aoi2222d1

.SUBCKT aoi2222d2 ZN  A1 A2 B1 B2 C1 C2 D1 D2 VDD VSS
MM24 VDD 2 4 VDD P l=0.18u w=1.09u 
MM23 4 3 VDD VDD P l=0.185937u w=1.152u 
MM22 VDD 4 ZN VDD P l=0.184173u w=1.984u 
MM21 VDD 4 ZN VDD P l=0.18u w=1.91u 
MM20 14 C2 3 VDD P l=0.185532u w=1.41u 
MM19 14 C1 3 VDD P l=0.18u w=1.34u 
MM18 14 D1 VDD VDD P l=0.184432u w=1.76u 
MM17 14 D2 VDD VDD P l=0.18u w=1.69u 
MM16 16 B2 VDD VDD P l=0.18u w=1.72u 
MM15 16 B1 VDD VDD P l=0.184358u w=1.79u 
MM14 16 A1 2 VDD P l=0.18u w=1.42u 
MM13 16 A2 2 VDD P l=0.185235u w=1.49u 
MM11 17 3 4 VSS N l=0.18u w=1.17u 
MM12 VSS 2 17 VSS N l=0.18u w=1.17u 
MM10 VSS 4 ZN VSS N l=0.18u w=1.19u 
MM9 VSS 4 ZN VSS N l=0.18u w=1.19u 
MM8 18 C2 VSS VSS N l=0.18u w=0.72u 
MM7 3 C1 18 VSS N l=0.18u w=0.72u 
MM6 3 D1 19 VSS N l=0.18u w=0.87u 
MM5 19 D2 VSS VSS N l=0.18u w=0.87u 
MM4 20 B2 VSS VSS N l=0.18u w=1u 
MM3 20 B1 2 VSS N l=0.186867u w=1.066u 
MM2 2 A1 21 VSS N l=0.18u w=0.72u 
MM1 VSS A2 21 VSS N l=0.18u w=0.72u 
.ENDS aoi2222d2

.SUBCKT aoi2222d4 ZN  A1 A2 B1 B2 C1 C2 D1 D2 VDD VSS
MM27 VDD 3 ZN VDD P l=0.184173u w=1.984u 
MM26 VDD 3 ZN VDD P l=0.18u w=1.91u 
MM25 VDD 3 ZN VDD P l=0.18u w=1.91u 
MM24 ZN 3 VDD VDD P l=0.184173u w=1.984u 
MM28 3 2 VDD VDD P l=0.18u w=1.09u 
MM23 VDD 4 3 VDD P l=0.185937u w=1.152u 
MM22 15 C2 4 VDD P l=0.185532u w=1.41u 
MM21 15 C1 4 VDD P l=0.18u w=1.34u 
MM20 VDD D1 15 VDD P l=0.184432u w=1.76u 
MM19 15 D2 VDD VDD P l=0.18u w=1.69u 
MM18 16 B2 VDD VDD P l=0.18u w=1.72u 
MM17 16 B1 VDD VDD P l=0.184358u w=1.79u 
MM16 16 A1 2 VDD P l=0.18u w=1.42u 
MM15 16 A2 2 VDD P l=0.185235u w=1.49u 
MM13 ZN 3 VSS VSS N l=0.187264u w=1.272u 
MM11 ZN 3 VSS VSS N l=0.18u w=1.19u 
MM12 VSS 3 ZN VSS N l=0.186551u w=1.264u 
MM10 ZN 3 VSS VSS N l=0.18u w=1.19u 
MM9 17 4 3 VSS N l=0.18u w=1.17u 
MM14 17 2 VSS VSS N l=0.18u w=1.17u 
MM8 18 C2 VSS VSS N l=0.18u w=0.72u 
MM7 18 C1 4 VSS N l=0.18u w=0.72u 
MM6 4 D1 19 VSS N l=0.18u w=0.87u 
MM5 VSS D2 19 VSS N l=0.18u w=0.87u 
MM4 20 B2 VSS VSS N l=0.18u w=1u 
MM3 20 B1 2 VSS N l=0.186867u w=1.066u 
MM2 2 A1 21 VSS N l=0.18u w=0.72u 
MM1 VSS A2 21 VSS N l=0.18u w=0.72u 
.ENDS aoi2222d4

.SUBCKT aoi222d1 ZN  A1 A2 B1 B2 C1 C2 VDD VSS
MM12 9 B2 10 VDD P l=0.18513u w=1.614u 
MM11 ZN A2 10 VDD P l=0.18u w=1.43u 
MM9 9 B1 10 VDD P l=0.18u w=1.54u 
MM10 ZN A1 10 VDD P l=0.1852u w=1.5u 
MM8 VDD C2 9 VDD P l=0.184043u w=1.692u 
MM7 VDD C1 9 VDD P l=0.187543u w=1.75u 
MM5 ZN C2 12 VSS N l=0.18u w=1.13u 
MM4 12 C1 VSS VSS N l=0.18u w=1.13u 
MM3 ZN A2 13 VSS N l=0.18u w=1.13u 
MM2 VSS A1 13 VSS N l=0.18u w=1.13u 
MM6 14 B2 VSS VSS N l=0.18u w=1.13u 
MM1 ZN B1 14 VSS N l=0.18u w=1.13u 
.ENDS aoi222d1

.SUBCKT aoi222d2 ZN  A1 A2 B1 B2 C1 C2 VDD VSS
MM18 10 C1 VDD VDD P l=0.18u w=1.71u 
MM16 10 B2 13 VDD P l=0.18513u w=1.614u 
MM17 10 C2 VDD VDD P l=0.184641u w=1.784u 
MM15 13 B1 10 VDD P l=0.18u w=1.54u 
MM14 7 6 VDD VDD P l=0.184483u w=1.74u 
MM13 VDD 7 ZN VDD P l=0.184483u w=1.74u 
MM12 VDD 7 ZN VDD P l=0.18u w=1.67u 
MM11 13 A1 6 VDD P l=0.18u w=1.48u 
MM10 13 A2 6 VDD P l=0.185032u w=1.55u 
MM9 14 C1 6 VSS N l=0.18u w=1.1u 
MM8 14 C2 VSS VSS N l=0.18u w=1.1u 
MM7 7 6 VSS VSS N l=0.18u w=1.54u 
MM6 VSS 7 ZN VSS N l=0.18u w=1.54u 
MM5 ZN 7 VSS VSS N l=0.18u w=1.54u 
MM4 6 A1 15 VSS N l=0.18u w=0.98u 
MM3 VSS A2 15 VSS N l=0.18u w=0.98u 
MM2 16 B2 VSS VSS N l=0.18u w=0.98u 
MM1 16 B1 6 VSS N l=0.18u w=0.98u 
.ENDS aoi222d2

.SUBCKT aoi222d4 ZN  A1 A2 B1 B2 C1 C2 VDD VSS
MM20 10 C2 VDD VDD P l=0.184641u w=1.784u 
MM19 10 C1 VDD VDD P l=0.18u w=1.71u 
MM18 10 B2 13 VDD P l=0.18513u w=1.614u 
MM17 13 B1 10 VDD P l=0.18u w=1.54u 
MM16 7 6 VDD VDD P l=0.184671u w=1.67u 
MM14 ZN 7 VDD VDD P l=0.183786u w=2.06u 
MM15 ZN 7 VDD VDD P l=0.183786u w=2.06u 
MM13 ZN 7 VDD VDD P l=0.18u w=1.99u 
MM12 13 A1 6 VDD P l=0.18u w=1.48u 
MM11 13 A2 6 VDD P l=0.185032u w=1.55u 
MM9 VSS 7 ZN VSS N l=0.18u w=1.61u 
MM8 VSS 7 ZN VSS N l=0.18u w=1.61u 
MM7 ZN 7 VSS VSS N l=0.18u w=1.61u 
MM10 14 C2 VSS VSS N l=0.18u w=1.1u 
MM6 14 C1 6 VSS N l=0.18u w=1.1u 
MM5 VSS 6 7 VSS N l=0.185417u w=1.44u 
MM4 6 A1 15 VSS N l=0.18u w=0.98u 
MM3 VSS A2 15 VSS N l=0.18u w=0.98u 
MM2 16 B2 VSS VSS N l=0.18u w=0.98u 
MM1 16 B1 6 VSS N l=0.18u w=0.98u 
.ENDS aoi222d4

.SUBCKT aoi22d1 ZN  A1 A2 B1 B2 VDD VSS
MM8 7 B2 VDD VDD P l=0.185132u w=1.52u 
MM7 7 B1 VDD VDD P l=0.184524u w=1.512u 
MM6 ZN A1 7 VDD P l=0.18u w=1.45u 
MM5 ZN A2 7 VDD P l=0.186796u w=1.545u 
MM4 9 B2 VSS VSS N l=0.188632u w=1.126u 
MM3 ZN B1 9 VSS N l=0.18u w=1.04u 
MM2 10 A1 ZN VSS N l=0.18u w=1.04u 
MM1 VSS A2 10 VSS N l=0.18u w=1.04u 
.ENDS aoi22d1

.SUBCKT aoi22d2 ZN  A1 A2 B1 B2 VDD VSS
MM14 8 A2 6 VDD P l=0.186796u w=1.545u 
MM13 6 A1 8 VDD P l=0.18u w=1.45u 
MM12 VDD B1 8 VDD P l=0.184524u w=1.512u 
MM11 VDD B2 8 VDD P l=0.185132u w=1.52u 
MM10 VDD 6 7 VDD P l=0.18u w=1.1u 
MM9 ZN 7 VDD VDD P l=0.183838u w=1.782u 
MM8 ZN 7 VDD VDD P l=0.183838u w=1.782u 
MM6 11 A1 6 VSS N l=0.18u w=1.04u 
MM5 6 B1 12 VSS N l=0.18u w=1.04u 
MM7 11 A2 VSS VSS N l=0.18u w=1.04u 
MM4 VSS B2 12 VSS N l=0.188632u w=1.126u 
MM3 VSS 6 7 VSS N l=0.18u w=0.88u 
MM2 VSS 7 ZN VSS N l=0.187013u w=1.386u 
MM1 VSS 7 ZN VSS N l=0.18u w=1.3u 
.ENDS aoi22d2

.SUBCKT aoi22d4 ZN  A1 A2 B1 B2 VDD VSS
MM16 VDD 2 3 VDD P l=0.18u w=1.45u 
MM15 VDD 3 ZN VDD P l=0.183786u w=2.06u 
MM14 ZN 3 VDD VDD P l=0.184459u w=2.072u 
MM13 ZN 3 VDD VDD P l=0.18u w=1.99u 
MM12 10 A2 2 VDD P l=0.186796u w=1.545u 
MM11 2 A1 10 VDD P l=0.18u w=1.45u 
MM10 VDD B1 10 VDD P l=0.184524u w=1.512u 
MM9 VDD B2 10 VDD P l=0.185132u w=1.52u 
MM8 3 2 VSS VSS N l=0.18u w=1.19u 
MM6 VSS 3 ZN VSS N l=0.184643u w=1.68u 
MM7 ZN 3 VSS VSS N l=0.185461u w=1.692u 
MM5 ZN 3 VSS VSS N l=0.18u w=1.61u 
MM3 11 A1 2 VSS N l=0.18u w=1.04u 
MM2 2 B1 12 VSS N l=0.18u w=1.04u 
MM4 11 A2 VSS VSS N l=0.18u w=1.04u 
MM1 VSS B2 12 VSS N l=0.188632u w=1.126u 
.ENDS aoi22d4

.SUBCKT aoi311d1 ZN  A B C1 C2 C3 VDD VSS
MM10 8 C1 VDD VDD P l=0.18u w=1.67u 
MM7 8 B 12 VDD P l=0.185235u w=1.49u 
MM9 VDD C3 8 VDD P l=0.184483u w=1.74u 
MM8 8 C2 VDD VDD P l=0.18u w=1.67u 
MM6 ZN A 12 VDD P l=0.185235u w=1.49u 
MM5 ZN C1 10 VSS N l=0.18u w=1.26u 
MM3 10 C2 11 VSS N l=0.185865u w=1.33u 
MM4 VSS C3 11 VSS N l=0.185865u w=1.33u 
MM2 VSS B ZN VSS N l=0.185865u w=1.33u 
MM1 VSS A ZN VSS N l=0.18u w=1.07u 
.ENDS aoi311d1

.SUBCKT aoi311d2 ZN  A B C1 C2 C3 VDD VSS
MM15 11 B 14 VDD P l=0.18u w=1.43u 
MM14 7 A 14 VDD P l=0.1852u w=1.5u 
MM16 VDD C3 11 VDD P l=0.18u w=1.63u 
MM13 VDD C2 11 VDD P l=0.184859u w=1.704u 
MM12 VDD C1 11 VDD P l=0.18u w=1.63u 
MM11 VDD 7 8 VDD P l=0.186096u w=1.122u 
MM10 ZN 8 VDD VDD P l=0.184216u w=1.85u 
MM9 VDD 8 ZN VDD P l=0.18u w=1.78u 
MM6 VSS A 7 VSS N l=0.18u w=0.98u 
MM8 VSS C3 12 VSS N l=0.18u w=1.04u 
MM5 13 C2 12 VSS N l=0.18u w=1.04u 
MM7 VSS B 7 VSS N l=0.187027u w=1.11u 
MM4 7 C1 13 VSS N l=0.18u w=1.04u 
MM3 8 7 VSS VSS N l=0.186446u w=1.21u 
MM2 VSS 8 ZN VSS N l=0.1852u w=1.5u 
MM1 ZN 8 VSS VSS N l=0.18u w=1.33u 
.ENDS aoi311d2

.SUBCKT aoi311d4 ZN  A B C1 C2 C3 VDD VSS
MM17 11 B 14 VDD P l=0.18u w=1.43u 
MM16 7 A 14 VDD P l=0.1852u w=1.5u 
MM18 VDD C3 11 VDD P l=0.18u w=1.63u 
MM15 11 C2 VDD VDD P l=0.184043u w=1.692u 
MM14 11 C1 VDD VDD P l=0.18u w=1.63u 
MM13 VDD 7 8 VDD P l=0.186096u w=1.122u 
MM12 ZN 8 VDD VDD P l=0.184236u w=2.068u 
MM11 VDD 8 ZN VDD P l=0.18u w=1.99u 
MM10 ZN 8 VDD VDD P l=0.18u w=1.99u 
MM7 VSS A 7 VSS N l=0.18u w=0.98u 
MM9 VSS C3 12 VSS N l=0.18u w=1.04u 
MM6 13 C2 12 VSS N l=0.18u w=1.04u 
MM8 VSS B 7 VSS N l=0.187027u w=1.11u 
MM5 7 C1 13 VSS N l=0.18u w=1.04u 
MM4 8 7 VSS VSS N l=0.186446u w=1.21u 
MM3 VSS 8 ZN VSS N l=0.18u w=1.41u 
MM2 VSS 8 ZN VSS N l=0.18527u w=1.48u 
MM1 ZN 8 VSS VSS N l=0.18u w=1.33u 
.ENDS aoi311d4

.SUBCKT aoi31d1 ZN  A B1 B2 B3 VDD VSS
MM8 6 B3 VDD VDD P l=0.18u w=1.15u 
MM7 6 B2 VDD VDD P l=0.185644u w=1.212u 
MM6 6 B1 VDD VDD P l=0.185644u w=1.212u 
MM5 ZN A 6 VDD P l=0.18u w=1.15u 
MM4 9 B3 VSS VSS N l=0.18u w=1.05u 
MM3 10 B2 9 VSS N l=0.18u w=1.05u 
MM2 10 B1 ZN VSS N l=0.18u w=1.05u 
MM1 ZN A VSS VSS N l=0.188163u w=1.132u 
.ENDS aoi31d1

.SUBCKT aoi31d2 ZN  A B1 B2 B3 VDD VSS
MM13 VDD 3 4 VDD P l=0.18u w=1.09u 
MM12 VDD 4 ZN VDD P l=0.185414u w=1.618u 
MM11 VDD 4 ZN VDD P l=0.18u w=1.54u 
MM14 10 B3 VDD VDD P l=0.18u w=1.15u 
MM10 10 B2 VDD VDD P l=0.185644u w=1.212u 
MM9 10 B1 VDD VDD P l=0.185644u w=1.212u 
MM8 3 A 10 VDD P l=0.18u w=1.15u 
MM6 VSS 3 4 VSS N l=0.18u w=0.91u 
MM5 ZN 4 VSS VSS N l=0.18602u w=1.216u 
MM4 ZN 4 VSS VSS N l=0.187424u w=0.986u 
MM7 VSS B3 11 VSS N l=0.18u w=1.11u 
MM3 11 B2 12 VSS N l=0.18u w=1.11u 
MM2 3 B1 12 VSS N l=0.18u w=1.11u 
MM1 3 A VSS VSS N l=0.187752u w=1.192u 
.ENDS aoi31d2

.SUBCKT aoi31d4 ZN  A B1 B2 B3 VDD VSS
MM16 VDD 2 3 VDD P l=0.18u w=1.09u 
MM15 ZN 3 VDD VDD P l=0.184012u w=2.064u 
MM14 ZN 3 VDD VDD P l=0.18u w=1.99u 
MM13 VDD 3 ZN VDD P l=0.183786u w=2.06u 
MM12 2 A 10 VDD P l=0.186393u w=1.22u 
MM11 VDD B1 10 VDD P l=0.18u w=1.15u 
MM10 10 B2 VDD VDD P l=0.18u w=1.15u 
MM9 VDD B3 10 VDD P l=0.186393u w=1.22u 
MM8 3 2 VSS VSS N l=0.18u w=0.91u 
MM6 VSS 3 ZN VSS N l=0.184643u w=1.68u 
MM7 ZN 3 VSS VSS N l=0.184917u w=1.684u 
MM5 ZN 3 VSS VSS N l=0.18u w=1.61u 
MM4 VSS A 2 VSS N l=0.186224u w=1.176u 
MM3 11 B1 2 VSS N l=0.18u w=1.11u 
MM2 12 B2 11 VSS N l=0.18u w=1.11u 
MM1 12 B3 VSS VSS N l=0.18u w=1.11u 
.ENDS aoi31d4

.SUBCKT aoi321d1 ZN  A B1 B2 C1 C2 C3 VDD VSS
MM12 VDD C1 9 VDD P l=0.185067u w=1.634u 
MM11 VDD C2 9 VDD P l=0.18u w=1.56u 
MM10 VDD C3 9 VDD P l=0.185067u w=1.634u 
MM9 9 B2 11 VDD P l=0.18u w=1.38u 
MM8 9 B1 11 VDD P l=0.185379u w=1.45u 
MM7 ZN A 11 VDD P l=0.185909u w=1.32u 
MM6 12 C1 ZN VSS N l=0.18u w=0.98u 
MM5 12 C2 13 VSS N l=0.18u w=0.98u 
MM4 13 C3 VSS VSS N l=0.18u w=0.98u 
MM3 ZN A VSS VSS N l=0.18u w=0.59u 
MM1 14 B1 ZN VSS N l=0.18u w=0.98u 
MM2 14 B2 VSS VSS N l=0.18u w=0.98u 
.ENDS aoi321d1

.SUBCKT aoi321d2 ZN  A B1 B2 C1 C2 C3 VDD VSS
MM18 VDD C2 10 VDD P l=0.18u w=1.56u 
MM17 VDD C1 10 VDD P l=0.185067u w=1.634u 
MM16 VDD C3 10 VDD P l=0.185067u w=1.634u 
MM15 10 B2 13 VDD P l=0.18u w=1.38u 
MM14 10 B1 13 VDD P l=0.185379u w=1.45u 
MM13 8 7 VDD VDD P l=0.185886u w=1.162u 
MM12 ZN 8 VDD VDD P l=0.18354u w=1.932u 
MM11 ZN 8 VDD VDD P l=0.18u w=1.87u 
MM10 7 A 13 VDD P l=0.185909u w=1.32u 
MM8 14 C1 7 VSS N l=0.18u w=0.98u 
MM9 14 C2 15 VSS N l=0.18u w=0.98u 
MM6 15 C3 VSS VSS N l=0.18u w=0.98u 
MM7 7 A VSS VSS N l=0.18u w=0.59u 
MM4 16 B1 7 VSS N l=0.18u w=0.98u 
MM5 16 B2 VSS VSS N l=0.18u w=0.98u 
MM3 VSS 7 8 VSS N l=0.186341u w=1.23u 
MM2 ZN 8 VSS VSS N l=0.185612u w=1.39u 
MM1 VSS 8 ZN VSS N l=0.18u w=1.32u 
.ENDS aoi321d2

.SUBCKT aoi321d4 ZN  A B1 B2 C1 C2 C3 VDD VSS
MM20 VDD C1 10 VDD P l=0.185067u w=1.634u 
MM19 VDD C2 10 VDD P l=0.18u w=1.56u 
MM18 VDD C3 10 VDD P l=0.185067u w=1.634u 
MM17 10 B2 13 VDD P l=0.18u w=1.38u 
MM16 10 B1 13 VDD P l=0.185379u w=1.45u 
MM15 8 7 VDD VDD P l=0.186667u w=1.17u 
MM14 ZN 8 VDD VDD P l=0.183786u w=2.06u 
MM13 VDD 8 ZN VDD P l=0.18u w=1.99u 
MM12 ZN 8 VDD VDD P l=0.183786u w=2.06u 
MM11 7 A 13 VDD P l=0.185909u w=1.32u 
MM10 14 C1 7 VSS N l=0.18u w=0.98u 
MM9 14 C2 15 VSS N l=0.18u w=0.98u 
MM7 15 C3 VSS VSS N l=0.18u w=0.98u 
MM8 7 A VSS VSS N l=0.18u w=0.59u 
MM5 16 B1 7 VSS N l=0.18u w=0.98u 
MM6 16 B2 VSS VSS N l=0.18u w=0.98u 
MM4 8 7 VSS VSS N l=0.185235u w=1.49u 
MM2 ZN 8 VSS VSS N l=0.184643u w=1.68u 
MM3 VSS 8 ZN VSS N l=0.184643u w=1.68u 
MM1 ZN 8 VSS VSS N l=0.18u w=1.61u 
.ENDS aoi321d4

.SUBCKT aoi322d1 ZN  A1 A2 B1 B2 C1 C2 C3 VDD VSS
MM13 VDD C1 10 VDD P l=0.18u w=1.65u 
MM12 10 C2 VDD VDD P l=0.184803u w=1.724u 
MM14 10 B2 11 VDD P l=0.185542u w=1.494u 
MM11 10 C3 VDD VDD P l=0.18u w=1.65u 
MM10 11 B1 10 VDD P l=0.18u w=1.42u 
MM9 ZN A1 11 VDD P l=0.18u w=1.52u 
MM8 ZN A2 11 VDD P l=0.184906u w=1.59u 
MM6 13 C1 ZN VSS N l=0.18u w=1.06u 
MM5 14 C2 13 VSS N l=0.18u w=1.06u 
MM4 14 C3 VSS VSS N l=0.18u w=1.06u 
MM3 ZN A1 15 VSS N l=0.18u w=0.82u 
MM2 VSS A2 15 VSS N l=0.18u w=0.82u 
MM1 ZN B1 16 VSS N l=0.18u w=1.06u 
MM7 16 B2 VSS VSS N l=0.18u w=1.06u 
.ENDS aoi322d1

.SUBCKT aoi322d2 ZN  A1 A2 B1 B2 C1 C2 C3 VDD VSS
MM20 11 C2 VDD VDD P l=0.184803u w=1.724u 
MM19 VDD C1 11 VDD P l=0.18u w=1.65u 
MM18 11 B2 14 VDD P l=0.185542u w=1.494u 
MM17 11 C3 VDD VDD P l=0.18u w=1.65u 
MM16 14 B1 11 VDD P l=0.18u w=1.42u 
MM15 VDD 7 8 VDD P l=0.186724u w=1.16u 
MM14 VDD 8 ZN VDD P l=0.185227u w=1.584u 
MM13 ZN 8 VDD VDD P l=0.18u w=1.51u 
MM12 14 A1 7 VDD P l=0.18u w=1.52u 
MM11 14 A2 7 VDD P l=0.184906u w=1.59u 
MM9 15 C1 7 VSS N l=0.18u w=1.06u 
MM10 16 C2 15 VSS N l=0.18u w=1.06u 
MM7 16 C3 VSS VSS N l=0.18u w=1.06u 
MM6 7 B1 17 VSS N l=0.18u w=1.06u 
MM5 7 A1 18 VSS N l=0.18u w=0.82u 
MM8 17 B2 VSS VSS N l=0.18u w=1.06u 
MM4 VSS A2 18 VSS N l=0.18u w=0.82u 
MM3 8 7 VSS VSS N l=0.18u w=1.05u 
MM2 VSS 8 ZN VSS N l=0.18u w=1.33u 
MM1 VSS 8 ZN VSS N l=0.18u w=1.33u 
.ENDS aoi322d2

.SUBCKT aoi322d4 ZN  A1 A2 B1 B2 C1 C2 C3 VDD VSS
MM22 11 C2 VDD VDD P l=0.184803u w=1.724u 
MM21 VDD C1 11 VDD P l=0.18u w=1.65u 
MM20 11 C3 VDD VDD P l=0.18u w=1.65u 
MM19 11 B2 14 VDD P l=0.185542u w=1.494u 
MM18 14 B1 11 VDD P l=0.18u w=1.42u 
MM17 VDD 7 8 VDD P l=0.186724u w=1.16u 
MM16 ZN 8 VDD VDD P l=0.184012u w=2.064u 
MM15 VDD 8 ZN VDD P l=0.18u w=1.99u 
MM14 VDD 8 ZN VDD P l=0.183786u w=2.06u 
MM13 7 A1 14 VDD P l=0.18u w=1.52u 
MM12 7 A2 14 VDD P l=0.184906u w=1.59u 
MM10 15 C1 7 VSS N l=0.18u w=1.06u 
MM11 17 C2 15 VSS N l=0.18u w=1.06u 
MM9 7 A1 16 VSS N l=0.18u w=0.82u 
MM8 VSS A2 16 VSS N l=0.18u w=0.82u 
MM7 17 C3 VSS VSS N l=0.18u w=1.06u 
MM5 7 B1 18 VSS N l=0.18u w=1.06u 
MM6 18 B2 VSS VSS N l=0.18u w=1.06u 
MM4 VSS 7 8 VSS N l=0.18u w=1.05u 
MM2 VSS 8 ZN VSS N l=0.184643u w=1.68u 
MM3 ZN 8 VSS VSS N l=0.184917u w=1.684u 
MM1 VSS 8 ZN VSS N l=0.18u w=1.61u 
.ENDS aoi322d4

.SUBCKT aoim211d1 ZN  A B C1 C2 VDD VSS
MM9 ZN A 9 VDD P l=0.188296u w=1.555u 
MM8 9 B 10 VDD P l=0.185166u w=1.51u 
MM10 VDD 2 10 VDD P l=0.185166u w=1.51u 
MM6 2 C1 11 VDD P l=0.185865u w=1.33u 
MM7 VDD C2 11 VDD P l=0.18u w=1.26u 
MM4 ZN A VSS VSS N l=0.187978u w=1.098u 
MM5 VSS 2 ZN VSS N l=0.18871u w=1.116u 
MM3 VSS B ZN VSS N l=0.18u w=1.03u 
MM2 2 C2 VSS VSS N l=0.18u w=1.13u 
MM1 2 C1 VSS VSS N l=0.1865u w=1.2u 
.ENDS aoim211d1

.SUBCKT aoim211d2 ZN  A B C1 C2 VDD VSS
MM16 7 A 11 VDD P l=0.188296u w=1.555u 
MM15 11 B 12 VDD P l=0.185166u w=1.51u 
MM14 VDD 4 12 VDD P l=0.185166u w=1.51u 
MM12 4 C1 13 VDD P l=0.185865u w=1.33u 
MM13 VDD C2 13 VDD P l=0.18u w=1.26u 
MM11 VDD 7 8 VDD P l=0.187222u w=1.08u 
MM10 ZN 8 VDD VDD P l=0.184815u w=1.62u 
MM9 ZN 8 VDD VDD P l=0.18u w=1.55u 
MM8 7 A VSS VSS N l=0.187978u w=1.098u 
MM7 7 B VSS VSS N l=0.18u w=1.04u 
MM6 7 4 VSS VSS N l=0.188632u w=1.126u 
MM5 VSS C2 4 VSS N l=0.18u w=1.13u 
MM4 VSS C1 4 VSS N l=0.1865u w=1.2u 
MM3 8 7 VSS VSS N l=0.18u w=0.91u 
MM2 ZN 8 VSS VSS N l=0.186993u w=1.184u 
MM1 ZN 8 VSS VSS N l=0.18u w=1.11u 
.ENDS aoim211d2

.SUBCKT aoim211d4 ZN  A B C1 C2 VDD VSS
MM18 7 A 11 VDD P l=0.188296u w=1.555u 
MM17 11 B 12 VDD P l=0.185166u w=1.51u 
MM16 VDD 4 12 VDD P l=0.185166u w=1.51u 
MM14 4 C1 13 VDD P l=0.185865u w=1.33u 
MM15 VDD C2 13 VDD P l=0.18u w=1.26u 
MM13 VDD 7 8 VDD P l=0.185u w=1.56u 
MM12 ZN 8 VDD VDD P l=0.183786u w=2.06u 
MM11 VDD 8 ZN VDD P l=0.18u w=1.99u 
MM10 ZN 8 VDD VDD P l=0.18u w=1.99u 
MM9 7 A VSS VSS N l=0.187978u w=1.098u 
MM8 7 B VSS VSS N l=0.18u w=1.03u 
MM7 7 4 VSS VSS N l=0.18871u w=1.116u 
MM6 VSS C2 4 VSS N l=0.18u w=1.13u 
MM5 VSS C1 4 VSS N l=0.1865u w=1.2u 
MM4 8 7 VSS VSS N l=0.18u w=1.09u 
MM2 ZN 8 VSS VSS N l=0.185778u w=1.35u 
MM3 VSS 8 ZN VSS N l=0.186115u w=1.354u 
MM1 ZN 8 VSS VSS N l=0.18u w=1.28u 
.ENDS aoim211d4

.SUBCKT aoim21d1 ZN  A B1 B2 VDD VSS
MM7 ZN A 8 VDD P l=0.18u w=1.54u 
MM8 8 2 VDD VDD P l=0.18u w=1.54u 
MM6 9 B2 VDD VDD P l=0.18u w=1.3u 
MM5 9 B1 2 VDD P l=0.185359u w=1.366u 
MM4 VSS 2 ZN VSS N l=0.187222u w=1.08u 
MM3 VSS A ZN VSS N l=0.18u w=1.01u 
MM2 VSS B2 2 VSS N l=0.18u w=1.09u 
MM1 VSS B1 2 VSS N l=0.186724u w=1.16u 
.ENDS aoim21d1

.SUBCKT aoim21d2 ZN  A B1 B2 VDD VSS
MM14 10 B2 VDD VDD P l=0.18u w=1.3u 
MM13 10 B1 5 VDD P l=0.185359u w=1.366u 
MM12 6 A 11 VDD P l=0.18u w=1.54u 
MM11 11 5 VDD VDD P l=0.18u w=1.54u 
MM10 7 6 VDD VDD P l=0.187222u w=1.08u 
MM9 VDD 7 ZN VDD P l=0.184815u w=1.62u 
MM8 ZN 7 VDD VDD P l=0.18u w=1.55u 
MM7 VSS B2 5 VSS N l=0.18u w=1.09u 
MM6 VSS B1 5 VSS N l=0.186724u w=1.16u 
MM5 VSS A 6 VSS N l=0.18u w=1.01u 
MM4 VSS 5 6 VSS N l=0.187222u w=1.08u 
MM3 7 6 VSS VSS N l=0.18u w=0.91u 
MM2 VSS 7 ZN VSS N l=0.186993u w=1.184u 
MM1 VSS 7 ZN VSS N l=0.18u w=1.11u 
.ENDS aoim21d2

.SUBCKT aoim21d4 ZN  A B1 B2 VDD VSS
MM16 3 2 VDD VDD P l=0.185u w=1.56u 
MM15 ZN 3 VDD VDD P l=0.183786u w=2.06u 
MM14 ZN 3 VDD VDD P l=0.18u w=1.99u 
MM13 VDD 3 ZN VDD P l=0.18u w=1.99u 
MM12 10 B2 VDD VDD P l=0.18u w=1.3u 
MM11 10 B1 7 VDD P l=0.185359u w=1.366u 
MM10 2 A 11 VDD P l=0.18u w=1.54u 
MM9 11 7 VDD VDD P l=0.18u w=1.54u 
MM8 3 2 VSS VSS N l=0.18u w=1.09u 
MM6 VSS 3 ZN VSS N l=0.185778u w=1.35u 
MM7 ZN 3 VSS VSS N l=0.186115u w=1.354u 
MM5 ZN 3 VSS VSS N l=0.18u w=1.28u 
MM4 VSS B2 7 VSS N l=0.18u w=1.09u 
MM3 VSS B1 7 VSS N l=0.186724u w=1.16u 
MM2 VSS A 2 VSS N l=0.18u w=1.01u 
MM1 VSS 7 2 VSS N l=0.187222u w=1.08u 
.ENDS aoim21d4

.SUBCKT aoim22d1 Z  A1 A2 B1 B2 VDD VSS
MM9 Z A2 9 VDD P l=0.184u w=1.95u 
MM8 Z A1 9 VDD P l=0.183522u w=1.942u 
MM10 VDD 2 9 VDD P l=0.184709u w=1.962u 
MM7 11 B2 VDD VDD P l=0.18u w=1.45u 
MM6 11 B1 2 VDD P l=0.18u w=1.45u 
MM5 Z 2 VSS VSS N l=0.18u w=1.13u 
MM3 10 A1 Z VSS N l=0.186168u w=1.576u 
MM4 10 A2 VSS VSS N l=0.185294u w=1.564u 
MM2 VSS B2 2 VSS N l=0.18u w=0.48u 
MM1 2 B1 VSS VSS N l=0.18u w=0.48u 
.ENDS aoim22d1

.SUBCKT aoim22d2 Z  A1 A2 B1 B2 VDD VSS
MM14 Z 3 VDD VDD P l=0.184815u w=1.62u 
MM13 Z 3 VDD VDD P l=0.18u w=1.55u 
MM15 3 B2 13 VDD P l=0.185455u w=1.43u 
MM12 VDD B1 13 VDD P l=0.185455u w=1.43u 
MM11 7 A2 VDD VDD P l=0.18u w=1.1u 
MM10 VDD A1 7 VDD P l=0.18u w=1.1u 
MM9 3 7 VDD VDD P l=0.185455u w=1.43u 
MM6 Z 3 VSS VSS N l=0.187374u w=1.188u 
MM5 VSS 3 Z VSS N l=0.18u w=1.11u 
MM7 VSS 7 10 VSS N l=0.18u w=1.23u 
MM4 3 B1 10 VSS N l=0.18u w=1.23u 
MM8 12 B2 3 VSS N l=0.18u w=1.23u 
MM3 VSS A2 11 VSS N l=0.18u w=0.96u 
MM2 7 A1 11 VSS N l=0.18u w=0.96u 
MM1 VSS 7 12 VSS N l=0.18u w=1.23u 
.ENDS aoim22d2

.SUBCKT aoim22d4 Z  A1 A2 B1 B2 VDD VSS
MM16 VDD 3 Z VDD P l=0.18356u w=2.056u 
MM15 VDD 3 Z VDD P l=0.18u w=1.99u 
MM14 VDD 3 Z VDD P l=0.18u w=1.99u 
MM13 7 A2 VDD VDD P l=0.18u w=1.1u 
MM12 VDD A1 7 VDD P l=0.18u w=1.1u 
MM17 VDD B1 13 VDD P l=0.185065u w=1.54u 
MM11 3 B2 13 VDD P l=0.185065u w=1.54u 
MM10 3 7 VDD VDD P l=0.185065u w=1.54u 
MM9 3 B1 10 VSS N l=0.18u w=1.23u 
MM8 VSS 7 10 VSS N l=0.18u w=1.23u 
MM7 Z 3 VSS VSS N l=0.185379u w=1.45u 
MM6 VSS 3 Z VSS N l=0.187043u w=1.312u 
MM5 Z 3 VSS VSS N l=0.18u w=1.38u 
MM4 11 A2 VSS VSS N l=0.18u w=0.95u 
MM3 7 A1 11 VSS N l=0.18u w=0.95u 
MM2 12 B2 3 VSS N l=0.18u w=1.23u 
MM1 VSS 7 12 VSS N l=0.18u w=1.23u 
.ENDS aoim22d4

.SUBCKT aoim2m11d1 ZN  A B C1 C2 VDD VSS
MM11 ZN A 10 VDD P l=0.18u w=1.52u 
MM10 11 4 10 VDD P l=0.18u w=1.52u 
MM9 11 5 VDD VDD P l=0.18u w=1.52u 
MM12 VDD C2 12 VDD P l=0.18552u w=1.326u 
MM8 5 C1 12 VDD P l=0.185865u w=1.33u 
MM7 4 B VDD VDD P l=0.185455u w=1.43u 
MM5 VSS A ZN VSS N l=0.186322u w=1.082u 
MM4 VSS 4 ZN VSS N l=0.18u w=1.02u 
MM3 VSS 5 ZN VSS N l=0.186322u w=1.082u 
MM6 5 C2 VSS VSS N l=0.18u w=0.98u 
MM2 5 C1 VSS VSS N l=0.18u w=0.98u 
MM1 4 B VSS VSS N l=0.18u w=0.98u 
.ENDS aoim2m11d1

.SUBCKT aoim2m11d2 ZN  A B C1 C2 VDD VSS
MM17 7 A 12 VDD P l=0.18u w=1.52u 
MM18 14 2 12 VDD P l=0.18u w=1.52u 
MM16 VDD C2 13 VDD P l=0.18552u w=1.326u 
MM15 6 C1 13 VDD P l=0.185865u w=1.33u 
MM14 14 6 VDD VDD P l=0.18u w=1.52u 
MM13 8 7 VDD VDD P l=0.187222u w=1.08u 
MM12 ZN 8 VDD VDD P l=0.184815u w=1.62u 
MM11 ZN 8 VDD VDD P l=0.18u w=1.55u 
MM10 2 B VDD VDD P l=0.185455u w=1.43u 
MM9 VSS 2 7 VSS N l=0.18u w=1.02u 
MM4 VSS 6 7 VSS N l=0.186322u w=1.082u 
MM8 VSS A 7 VSS N l=0.186322u w=1.082u 
MM7 6 C2 VSS VSS N l=0.18u w=0.98u 
MM6 6 C1 VSS VSS N l=0.18u w=0.98u 
MM5 2 B VSS VSS N l=0.18u w=0.98u 
MM3 8 7 VSS VSS N l=0.18u w=0.83u 
MM2 ZN 8 VSS VSS N l=0.186993u w=1.184u 
MM1 ZN 8 VSS VSS N l=0.18u w=1.11u 
.ENDS aoim2m11d2

.SUBCKT aoim2m11d4 ZN  A B C1 C2 VDD VSS
MM20 7 A 13 VDD P l=0.18u w=1.52u 
MM19 VDD C2 12 VDD P l=0.18552u w=1.326u 
MM18 6 C1 12 VDD P l=0.185865u w=1.33u 
MM17 14 5 13 VDD P l=0.18u w=1.52u 
MM16 14 6 VDD VDD P l=0.18u w=1.52u 
MM15 8 7 VDD VDD P l=0.18629u w=1.24u 
MM14 VDD 8 ZN VDD P l=0.183786u w=2.06u 
MM13 ZN 8 VDD VDD P l=0.18u w=1.99u 
MM12 ZN 8 VDD VDD P l=0.18u w=1.99u 
MM11 5 B VDD VDD P l=0.185455u w=1.43u 
MM10 VSS A 7 VSS N l=0.186322u w=1.082u 
MM9 6 C2 VSS VSS N l=0.18u w=0.98u 
MM8 6 C1 VSS VSS N l=0.18u w=0.98u 
MM7 5 B VSS VSS N l=0.18u w=0.98u 
MM6 VSS 5 7 VSS N l=0.18u w=1.02u 
MM5 VSS 6 7 VSS N l=0.186322u w=1.082u 
MM4 8 7 VSS VSS N l=0.18u w=0.83u 
MM2 ZN 8 VSS VSS N l=0.185652u w=1.38u 
MM3 ZN 8 VSS VSS N l=0.185983u w=1.384u 
MM1 VSS 8 ZN VSS N l=0.18u w=1.31u 
.ENDS aoim2m11d4

.SUBCKT aoim311d1 ZN  A B C1 C2 C3 VDD VSS
MM11 ZN A 10 VDD P l=0.18u w=1.97u 
MM10 11 B 10 VDD P l=0.18u w=1.97u 
MM12 11 2 VDD VDD P l=0.18u w=1.97u 
MM9 12 C3 VDD VDD P l=0.18u w=1.36u 
MM8 13 C2 12 VDD P l=0.18u w=1.36u 
MM7 13 C1 2 VDD P l=0.18u w=1.36u 
MM6 VSS 2 ZN VSS N l=0.186278u w=1.166u 
MM5 ZN A VSS VSS N l=0.186278u w=1.166u 
MM4 ZN B VSS VSS N l=0.18u w=1.1u 
MM3 VSS C3 2 VSS N l=0.18u w=0.8u 
MM2 VSS C2 2 VSS N l=0.18u w=1.18u 
MM1 VSS C1 2 VSS N l=0.186724u w=1.16u 
.ENDS aoim311d1

.SUBCKT aoim311d2 ZN  A B C1 C2 C3 VDD VSS
MM17 12 A 8 VDD P l=0.18u w=1.24u 
MM18 13 B 12 VDD P l=0.18u w=1.24u 
MM16 13 4 VDD VDD P l=0.18u w=1.24u 
MM15 VDD C3 14 VDD P l=0.18u w=1.24u 
MM14 15 C2 14 VDD P l=0.18u w=1.24u 
MM13 15 C1 4 VDD P l=0.18u w=1.24u 
MM12 9 8 VDD VDD P l=0.185011u w=1.748u 
MM11 ZN 9 VDD VDD P l=0.184875u w=1.6u 
MM10 ZN 9 VDD VDD P l=0.18u w=1.67u 
MM9 8 B VSS VSS N l=0.186254u w=1.324u 
MM8 8 A VSS VSS N l=0.18u w=1.25u 
MM7 VSS 8 9 VSS N l=0.185562u w=1.316u 
MM6 ZN 9 VSS VSS N l=0.186254u w=1.324u 
MM5 VSS 9 ZN VSS N l=0.18u w=1.25u 
MM4 VSS 4 8 VSS N l=0.18u w=1.14u 
MM3 VSS C3 4 VSS N l=0.18u w=0.98u 
MM2 VSS C2 4 VSS N l=0.18u w=1.08u 
MM1 VSS C1 4 VSS N l=0.186387u w=1.146u 
.ENDS aoim311d2

.SUBCKT aoim311d4 ZN  A B C1 C2 C3 VDD VSS
MM20 14 A 8 VDD P l=0.186746u w=1.841u 
MM19 12 C3 VDD VDD P l=0.18u w=1.29u 
MM18 12 C2 13 VDD P l=0.18u w=1.29u 
MM17 7 C1 13 VDD P l=0.185735u w=1.36u 
MM16 15 B 14 VDD P l=0.18u w=1.83u 
MM15 15 7 VDD VDD P l=0.18u w=1.83u 
MM14 VDD 8 9 VDD P l=0.187535u w=2.134u 
MM13 ZN 9 VDD VDD P l=0.185256u w=2.089u 
MM12 VDD 9 ZN VDD P l=0.18u w=1.99u 
MM11 VDD 9 ZN VDD P l=0.186471u w=2.114u 
MM10 VSS A 8 VSS N l=0.18629u w=1.24u 
MM9 VSS C3 7 VSS N l=0.18u w=1.08u 
MM8 7 C2 VSS VSS N l=0.187175u w=1.154u 
MM7 7 C1 VSS VSS N l=0.18u w=1.08u 
MM6 VSS B 8 VSS N l=0.18u w=1.17u 
MM5 8 7 VSS VSS N l=0.18629u w=1.24u 
MM4 9 8 VSS VSS N l=0.185571u w=1.4u 
MM2 VSS 9 ZN VSS N l=0.18u w=1.33u 
MM3 VSS 9 ZN VSS N l=0.185244u w=1.396u 
MM1 ZN 9 VSS VSS N l=0.18u w=1.33u 
.ENDS aoim311d4

.SUBCKT aoim31d1 ZN  A B1 B2 B3 VDD VSS
MM9 ZN A 9 VDD P l=0.184465u w=1.532u 
MM8 9 4 VDD VDD P l=0.18u w=1.47u 
MM10 10 B3 VDD VDD P l=0.184494u w=1.522u 
MM7 10 B2 11 VDD P l=0.18u w=1.46u 
MM6 4 B1 11 VDD P l=0.184494u w=1.522u 
MM4 VSS A ZN VSS N l=0.185787u w=1.182u 
MM3 ZN 4 VSS VSS N l=0.18u w=1.12u 
MM5 4 B3 VSS VSS N l=0.186172u w=1.186u 
MM2 4 B2 VSS VSS N l=0.18u w=1.12u 
MM1 4 B1 VSS VSS N l=0.186555u w=1.19u 
.ENDS aoim31d1

.SUBCKT aoim31d2 ZN  A B1 B2 B3 VDD VSS
MM16 7 A 13 VDD P l=0.184465u w=1.532u 
MM15 11 B3 VDD VDD P l=0.184494u w=1.522u 
MM14 11 B2 12 VDD P l=0.18u w=1.46u 
MM13 6 B1 12 VDD P l=0.184494u w=1.522u 
MM12 13 6 VDD VDD P l=0.18u w=1.47u 
MM11 VDD 7 8 VDD P l=0.187222u w=1.08u 
MM10 ZN 8 VDD VDD P l=0.184815u w=1.62u 
MM9 ZN 8 VDD VDD P l=0.18u w=1.55u 
MM7 6 B3 VSS VSS N l=0.186172u w=1.186u 
MM6 6 B2 VSS VSS N l=0.18u w=1.12u 
MM5 6 B1 VSS VSS N l=0.186555u w=1.19u 
MM8 VSS A 7 VSS N l=0.185787u w=1.182u 
MM4 7 6 VSS VSS N l=0.18u w=1.12u 
MM3 8 7 VSS VSS N l=0.18u w=0.91u 
MM2 ZN 8 VSS VSS N l=0.186993u w=1.184u 
MM1 ZN 8 VSS VSS N l=0.18u w=1.11u 
.ENDS aoim31d2

.SUBCKT aoim31d4 ZN  A B1 B2 B3 VDD VSS
MM18 11 B3 VDD VDD P l=0.184494u w=1.522u 
MM17 11 B2 12 VDD P l=0.18u w=1.46u 
MM16 6 B1 12 VDD P l=0.184494u w=1.522u 
MM15 7 A 13 VDD P l=0.184465u w=1.532u 
MM14 13 6 VDD VDD P l=0.18u w=1.47u 
MM13 VDD 7 8 VDD P l=0.18661u w=1.18u 
MM12 ZN 8 VDD VDD P l=0.183786u w=2.06u 
MM11 VDD 8 ZN VDD P l=0.18u w=1.99u 
MM10 ZN 8 VDD VDD P l=0.18u w=1.99u 
MM9 6 B3 VSS VSS N l=0.186172u w=1.186u 
MM8 6 B2 VSS VSS N l=0.18u w=1.12u 
MM7 6 B1 VSS VSS N l=0.186555u w=1.19u 
MM6 VSS A 7 VSS N l=0.185787u w=1.182u 
MM5 7 6 VSS VSS N l=0.18u w=1.12u 
MM4 8 7 VSS VSS N l=0.18u w=0.83u 
MM2 ZN 8 VSS VSS N l=0.185778u w=1.35u 
MM3 VSS 8 ZN VSS N l=0.186115u w=1.354u 
MM1 ZN 8 VSS VSS N l=0.18u w=1.28u 
.ENDS aoim31d4

.SUBCKT aoim3m11d1 ZN  A B C1 C2 C3 VDD VSS
MM13 ZN A 11 VDD P l=0.18u w=1.81u 
MM12 11 4 12 VDD P l=0.186839u w=1.93u 
MM11 VDD 5 12 VDD P l=0.187073u w=1.934u 
MM14 VDD C3 13 VDD P l=0.18u w=1.66u 
MM10 14 C2 13 VDD P l=0.18u w=1.66u 
MM9 14 C1 5 VDD P l=0.18u w=1.66u 
MM8 4 B VDD VDD P l=0.18u w=1.11u 
MM7 VSS C3 5 VSS N l=0.18u w=0.79u 
MM6 4 B VSS VSS N l=0.186387u w=1.146u 
MM5 5 C2 VSS VSS N l=0.187565u w=1.158u 
MM4 5 C1 VSS VSS N l=0.18u w=1.08u 
MM3 VSS A ZN VSS N l=0.186501u w=1.126u 
MM2 VSS 4 ZN VSS N l=0.186501u w=1.126u 
MM1 ZN 5 VSS VSS N l=0.18u w=1.06u 
.ENDS aoim3m11d1

.SUBCKT aoim3m11d2 ZN  A B C1 C2 C3 VDD VSS
MM20 13 2 14 VDD P l=0.187539u w=1.942u 
MM19 8 A 13 VDD P l=0.184884u w=1.892u 
MM18 VDD 4 14 VDD P l=0.188u w=1.95u 
MM17 15 C3 VDD VDD P l=0.18u w=1.66u 
MM16 16 C2 15 VDD P l=0.18u w=1.66u 
MM15 16 C1 4 VDD P l=0.18u w=1.66u 
MM14 VDD 8 9 VDD P l=0.1865u w=1.2u 
MM13 ZN 9 VDD VDD P l=0.184815u w=1.62u 
MM12 VDD 9 ZN VDD P l=0.18u w=1.55u 
MM11 2 B VDD VDD P l=0.18u w=1.11u 
MM9 VSS 8 9 VSS N l=0.18u w=0.91u 
MM8 VSS 9 ZN VSS N l=0.186993u w=1.184u 
MM7 VSS 9 ZN VSS N l=0.18u w=1.11u 
MM10 VSS 2 8 VSS N l=0.186501u w=1.126u 
MM6 VSS A 8 VSS N l=0.186501u w=1.126u 
MM5 8 4 VSS VSS N l=0.18u w=1.06u 
MM4 2 B VSS VSS N l=0.186387u w=1.146u 
MM3 VSS C3 4 VSS N l=0.18u w=0.79u 
MM2 4 C2 VSS VSS N l=0.187565u w=1.158u 
MM1 4 C1 VSS VSS N l=0.18u w=1.08u 
.ENDS aoim3m11d2

.SUBCKT aoim3m11d4 ZN  A B C1 C2 C3 VDD VSS
MM22 13 A 8 VDD P l=0.183654u w=1.872u 
MM21 13 3 14 VDD P l=0.187539u w=1.942u 
MM20 VDD 4 14 VDD P l=0.18777u w=1.946u 
MM19 15 C3 VDD VDD P l=0.18u w=1.66u 
MM18 16 C2 15 VDD P l=0.18u w=1.66u 
MM17 16 C1 4 VDD P l=0.18u w=1.66u 
MM16 9 8 VDD VDD P l=0.18629u w=1.24u 
MM15 ZN 9 VDD VDD P l=0.183786u w=2.06u 
MM14 ZN 9 VDD VDD P l=0.18u w=1.99u 
MM13 VDD 9 ZN VDD P l=0.18u w=1.99u 
MM12 3 B VDD VDD P l=0.18u w=1.11u 
MM11 VSS A 8 VSS N l=0.186501u w=1.126u 
MM10 VSS 3 8 VSS N l=0.186501u w=1.126u 
MM9 8 4 VSS VSS N l=0.18u w=1.06u 
MM8 9 8 VSS VSS N l=0.18u w=0.99u 
MM6 VSS 9 ZN VSS N l=0.185778u w=1.35u 
MM7 ZN 9 VSS VSS N l=0.186115u w=1.354u 
MM5 ZN 9 VSS VSS N l=0.18u w=1.28u 
MM4 3 B VSS VSS N l=0.186387u w=1.146u 
MM3 VSS C3 4 VSS N l=0.18u w=0.79u 
MM2 4 C2 VSS VSS N l=0.187565u w=1.158u 
MM1 4 C1 VSS VSS N l=0.18u w=1.08u 
.ENDS aoim3m11d4

.SUBCKT aon211d1 ZN  A B C1 C2 VDD VSS
MM8 VDD A ZN VDD P l=0.184968u w=1.57u 
MM7 ZN B 6 VDD P l=0.18u w=1.5u 
MM6 VDD C2 6 VDD P l=0.18526u w=1.574u 
MM5 VDD C1 6 VDD P l=0.184968u w=1.57u 
MM1 8 C1 10 VSS N l=0.188868u w=1.042u 
MM4 ZN A 8 VSS N l=0.186264u w=1.092u 
MM3 VSS B 8 VSS N l=0.186264u w=1.092u 
MM2 VSS C2 10 VSS N l=0.18u w=0.96u 
.ENDS aon211d1

.SUBCKT aon211d2 ZN  A B C1 C2 VDD VSS
MM14 VDD A 6 VDD P l=0.184968u w=1.57u 
MM13 6 B 11 VDD P l=0.18u w=1.5u 
MM12 VDD C2 11 VDD P l=0.18526u w=1.574u 
MM11 VDD C1 11 VDD P l=0.184968u w=1.57u 
MM10 7 6 VDD VDD P l=0.185886u w=1.162u 
MM9 ZN 7 VDD VDD P l=0.183838u w=1.782u 
MM8 ZN 7 VDD VDD P l=0.183838u w=1.782u 
MM4 10 C1 12 VSS N l=0.188235u w=1.122u 
MM7 6 A 10 VSS N l=0.186441u w=1.062u 
MM6 VSS B 10 VSS N l=0.186441u w=1.062u 
MM5 VSS C2 12 VSS N l=0.18u w=1.04u 
MM3 7 6 VSS VSS N l=0.18u w=0.88u 
MM2 ZN 7 VSS VSS N l=0.187386u w=1.316u 
MM1 ZN 7 VSS VSS N l=0.18u w=1.23u 
.ENDS aon211d2

.SUBCKT aon211d4 ZN  A B C1 C2 VDD VSS
MM16 3 2 VDD VDD P l=0.185886u w=1.162u 
MM15 ZN 3 VDD VDD P l=0.183333u w=2.052u 
MM14 ZN 3 VDD VDD P l=0.18u w=1.99u 
MM13 VDD 3 ZN VDD P l=0.184012u w=2.064u 
MM12 VDD A 2 VDD P l=0.18526u w=1.574u 
MM11 2 B 11 VDD P l=0.18u w=1.5u 
MM10 VDD C2 11 VDD P l=0.184968u w=1.57u 
MM9 VDD C1 11 VDD P l=0.184968u w=1.57u 
MM8 3 2 VSS VSS N l=0.18u w=0.88u 
MM6 VSS 3 ZN VSS N l=0.185983u w=1.384u 
MM7 ZN 3 VSS VSS N l=0.186963u w=1.396u 
MM5 ZN 3 VSS VSS N l=0.18u w=1.31u 
MM1 10 C1 12 VSS N l=0.188235u w=1.122u 
MM4 2 A 10 VSS N l=0.186441u w=1.062u 
MM3 VSS B 10 VSS N l=0.186441u w=1.062u 
MM2 VSS C2 12 VSS N l=0.18u w=1.04u 
.ENDS aon211d4

.SUBCKT aor211d1 Z  A B C1 C2 VDD VSS
MM9 7 C2 VDD VDD P l=0.185652u w=1.38u 
MM10 7 C1 VDD VDD P l=0.18u w=1.34u 
MM8 11 B 7 VDD P l=0.184671u w=1.67u 
MM7 11 A 6 VDD P l=0.184671u w=1.67u 
MM6 VDD 6 Z VDD P l=0.185417u w=1.44u 
MM5 10 C1 6 VSS N l=0.18u w=1.04u 
MM4 10 C2 VSS VSS N l=0.18u w=1.04u 
MM3 Z 6 VSS VSS N l=0.18u w=0.94u 
MM2 6 B VSS VSS N l=0.18u w=1.04u 
MM1 6 A VSS VSS N l=0.187222u w=1.08u 
.ENDS aor211d1

.SUBCKT aor211d2 Z  A B C1 C2 VDD VSS
MM12 7 C2 VDD VDD P l=0.186867u w=1.3325u 
MM11 VDD 3 Z VDD P l=0.184875u w=1.6u 
MM10 VDD 3 Z VDD P l=0.18u w=1.53u 
MM9 7 C1 VDD VDD P l=0.18u w=1.21u 
MM8 11 B 7 VDD P l=0.184815u w=1.62u 
MM7 11 A 3 VDD P l=0.184815u w=1.62u 
MM5 Z 3 VSS VSS N l=0.18u w=0.99u 
MM4 Z 3 VSS VSS N l=0.18u w=0.99u 
MM6 10 C2 VSS VSS N l=0.18u w=1.11u 
MM3 3 C1 10 VSS N l=0.18u w=1.11u 
MM2 3 B VSS VSS N l=0.18u w=1.11u 
MM1 3 A VSS VSS N l=0.185886u w=1.162u 
.ENDS aor211d2

.SUBCKT aor211d4 Z  A B C1 C2 VDD VSS
MM14 7 C2 VDD VDD P l=0.186047u w=1.29u 
MM13 VDD C1 7 VDD P l=0.187687u w=1.202u 
MM12 11 B 7 VDD P l=0.18u w=1.6u 
MM11 11 A 6 VDD P l=0.18u w=1.6u 
MM10 VDD 6 Z VDD P l=0.184682u w=2.076u 
MM9 Z 6 VDD VDD P l=0.18u w=1.99u 
MM8 VDD 6 Z VDD P l=0.18u w=1.99u 
MM6 Z 6 VSS VSS N l=0.185571u w=1.4u 
MM5 Z 6 VSS VSS N l=0.18u w=1.33u 
MM4 Z 6 VSS VSS N l=0.18u w=1.33u 
MM7 VSS C2 10 VSS N l=0.18u w=1.05u 
MM3 10 C1 6 VSS N l=0.18u w=1.05u 
MM2 VSS B 6 VSS N l=0.18u w=1.05u 
MM1 VSS A 6 VSS N l=0.186964u w=1.12u 
.ENDS aor211d4

.SUBCKT aor21d1 Z  A B1 B2 VDD VSS
MM8 VDD B2 6 VDD P l=0.18624u w=1.25u 
MM7 6 B1 VDD VDD P l=0.18u w=1.18u 
MM6 6 A 5 VDD P l=0.185875u w=1.246u 
MM5 VDD 5 Z VDD P l=0.185235u w=1.49u 
MM3 Z 5 VSS VSS N l=0.18u w=0.97u 
MM4 9 B2 VSS VSS N l=0.18u w=1.04u 
MM2 9 B1 5 VSS N l=0.18u w=1.04u 
MM1 VSS A 5 VSS N l=0.186207u w=1.102u 
.ENDS aor21d1

.SUBCKT aor21d2 Z  A B1 B2 VDD VSS
MM10 VDD B2 6 VDD P l=0.18624u w=1.25u 
MM9 6 B1 VDD VDD P l=0.18u w=1.18u 
MM8 6 A 5 VDD P l=0.185875u w=1.246u 
MM7 Z 5 VDD VDD P l=0.185235u w=1.49u 
MM6 VDD 5 Z VDD P l=0.18u w=1.42u 
MM4 VSS 5 Z VSS N l=0.18u w=0.97u 
MM3 VSS 5 Z VSS N l=0.18u w=0.97u 
MM5 9 B2 VSS VSS N l=0.18u w=1.04u 
MM2 9 B1 5 VSS N l=0.18u w=1.04u 
MM1 VSS A 5 VSS N l=0.186207u w=1.102u 
.ENDS aor21d2

.SUBCKT aor21d4 Z  A B1 B2 VDD VSS
MM12 6 B2 VDD VDD P l=0.186094u w=1.28u 
MM11 6 B1 VDD VDD P l=0.187152u w=1.292u 
MM10 5 A 6 VDD P l=0.18u w=1.21u 
MM9 VDD 5 Z VDD P l=0.184682u w=2.076u 
MM8 VDD 5 Z VDD P l=0.18u w=1.99u 
MM7 Z 5 VDD VDD P l=0.18u w=1.99u 
MM5 VSS 5 Z VSS N l=0.185571u w=1.4u 
MM4 Z 5 VSS VSS N l=0.18u w=1.33u 
MM3 Z 5 VSS VSS N l=0.18u w=1.33u 
MM6 9 B2 VSS VSS N l=0.18u w=1u 
MM2 9 B1 5 VSS N l=0.18u w=1u 
MM1 VSS A 5 VSS N l=0.18u w=1u 
.ENDS aor21d4

.SUBCKT aor221d1 Z  A B1 B2 C1 C2 VDD VSS
MM12 Z 2 VDD VDD P l=0.184937u w=1.58u 
MM11 8 C2 VDD VDD P l=0.18u w=1.56u 
MM10 VDD C1 8 VDD P l=0.184785u w=1.63u 
MM9 2 A 11 VDD P l=0.184893u w=1.496u 
MM8 8 B2 11 VDD P l=0.184785u w=1.63u 
MM7 8 B1 11 VDD P l=0.18u w=1.56u 
MM6 VSS 2 Z VSS N l=0.187222u w=1.08u 
MM5 VSS C2 12 VSS N l=0.18u w=1.01u 
MM4 12 C1 2 VSS N l=0.18u w=1.01u 
MM2 VSS B2 13 VSS N l=0.18u w=0.91u 
MM1 2 B1 13 VSS N l=0.18u w=0.91u 
MM3 2 A VSS VSS N l=0.18u w=0.91u 
.ENDS aor221d1

.SUBCKT aor221d2 Z  A B1 B2 C1 C2 VDD VSS
MM13 Z 3 VDD VDD P l=0.184243u w=1.612u 
MM12 Z 3 VDD VDD P l=0.184815u w=1.62u 
MM14 VDD C1 8 VDD P l=0.184785u w=1.63u 
MM11 8 C2 VDD VDD P l=0.18u w=1.56u 
MM10 3 A 11 VDD P l=0.184893u w=1.496u 
MM9 8 B2 11 VDD P l=0.184785u w=1.63u 
MM8 8 B1 11 VDD P l=0.18u w=1.56u 
MM7 12 C1 3 VSS N l=0.18u w=1.01u 
MM6 VSS 3 Z VSS N l=0.187638u w=1.084u 
MM5 VSS 3 Z VSS N l=0.187222u w=1.08u 
MM4 VSS C2 12 VSS N l=0.18u w=1.01u 
MM2 VSS B2 13 VSS N l=0.18u w=0.91u 
MM1 3 B1 13 VSS N l=0.18u w=0.91u 
MM3 3 A VSS VSS N l=0.18u w=0.91u 
.ENDS aor221d2

.SUBCKT aor221d4 Z  A B1 B2 C1 C2 VDD VSS
MM16 8 C1 VDD VDD P l=0.184785u w=1.63u 
MM15 8 C2 VDD VDD P l=0.18u w=1.56u 
MM14 Z 4 VDD VDD P l=0.183333u w=2.052u 
MM13 Z 4 VDD VDD P l=0.18u w=1.99u 
MM12 VDD 4 Z VDD P l=0.183786u w=2.06u 
MM11 11 A 4 VDD P l=0.184893u w=1.496u 
MM10 11 B1 8 VDD P l=0.18u w=1.56u 
MM9 8 B2 11 VDD P l=0.184785u w=1.63u 
MM8 12 C1 4 VSS N l=0.18u w=1.01u 
MM7 VSS C2 12 VSS N l=0.18u w=1.01u 
MM5 VSS 4 Z VSS N l=0.185612u w=1.39u 
MM6 VSS 4 Z VSS N l=0.185281u w=1.386u 
MM4 Z 4 VSS VSS N l=0.184949u w=1.382u 
MM3 4 A VSS VSS N l=0.18u w=0.91u 
MM2 4 B1 13 VSS N l=0.18u w=0.91u 
MM1 VSS B2 13 VSS N l=0.18u w=0.91u 
.ENDS aor221d4

.SUBCKT aor222d1 Z  A1 A2 B1 B2 C1 C2 VDD VSS
MM13 9 C2 VDD VDD P l=0.18u w=1.52u 
MM14 12 B2 9 VDD P l=0.18u w=1.52u 
MM12 9 C1 VDD VDD P l=0.185194u w=1.594u 
MM11 12 B1 9 VDD P l=0.184906u w=1.59u 
MM10 VDD 6 Z VDD P l=0.185098u w=1.53u 
MM9 6 A1 12 VDD P l=0.18u w=1.41u 
MM8 6 A2 12 VDD P l=0.18527u w=1.48u 
MM6 6 A1 13 VSS N l=0.18u w=0.86u 
MM5 VSS A2 13 VSS N l=0.18u w=0.86u 
MM7 14 B2 VSS VSS N l=0.18u w=0.86u 
MM4 14 B1 6 VSS N l=0.18u w=0.86u 
MM3 Z 6 VSS VSS N l=0.18u w=0.96u 
MM2 15 C2 VSS VSS N l=0.18u w=0.96u 
MM1 6 C1 15 VSS N l=0.18u w=0.96u 
.ENDS aor222d1

.SUBCKT aor222d2 Z  A1 A2 B1 B2 C1 C2 VDD VSS
MM16 9 C2 VDD VDD P l=0.18u w=1.52u 
MM15 9 C1 VDD VDD P l=0.185194u w=1.594u 
MM14 12 B2 9 VDD P l=0.18u w=1.52u 
MM13 12 B1 9 VDD P l=0.184906u w=1.59u 
MM12 VDD 6 Z VDD P l=0.185098u w=1.53u 
MM11 VDD 6 Z VDD P l=0.18u w=1.46u 
MM10 6 A1 12 VDD P l=0.18u w=1.41u 
MM9 6 A2 12 VDD P l=0.18527u w=1.48u 
MM8 Z 6 VSS VSS N l=0.18u w=0.96u 
MM7 Z 6 VSS VSS N l=0.18u w=0.96u 
MM6 13 C2 VSS VSS N l=0.18u w=0.96u 
MM5 6 C1 13 VSS N l=0.18u w=0.96u 
MM4 6 A1 14 VSS N l=0.18u w=0.86u 
MM3 VSS A2 14 VSS N l=0.18u w=0.86u 
MM2 15 B2 VSS VSS N l=0.18u w=0.86u 
MM1 15 B1 6 VSS N l=0.18u w=0.86u 
.ENDS aor222d2

.SUBCKT aor222d4 Z  A1 A2 B1 B2 C1 C2 VDD VSS
MM17 9 C2 VDD VDD P l=0.18u w=1.45u 
MM18 9 C1 VDD VDD P l=0.185433u w=1.524u 
MM16 12 B2 9 VDD P l=0.18u w=1.45u 
MM15 12 B1 9 VDD P l=0.185132u w=1.52u 
MM14 VDD 6 Z VDD P l=0.184012u w=2.064u 
MM13 VDD 6 Z VDD P l=0.18u w=1.99u 
MM12 VDD 6 Z VDD P l=0.183786u w=2.06u 
MM11 6 A1 12 VDD P l=0.18u w=1.41u 
MM10 6 A2 12 VDD P l=0.18527u w=1.48u 
MM9 6 C1 13 VSS N l=0.18u w=1.61u 
MM8 VSS C2 13 VSS N l=0.18u w=1.61u 
MM7 VSS 6 Z VSS N l=0.184643u w=1.68u 
MM6 VSS 6 Z VSS N l=0.18u w=1.61u 
MM5 VSS 6 Z VSS N l=0.18u w=1.61u 
MM4 6 A1 14 VSS N l=0.18u w=0.86u 
MM3 VSS A2 14 VSS N l=0.18u w=0.86u 
MM2 15 B2 VSS VSS N l=0.18u w=0.86u 
MM1 15 B1 6 VSS N l=0.18u w=0.86u 
.ENDS aor222d4

.SUBCKT aor22d1 Z  A1 A2 B1 B2 VDD VSS
MM10 7 A2 6 VDD P l=0.18u w=1.35u 
MM9 7 A1 6 VDD P l=0.185815u w=1.424u 
MM8 VDD B1 7 VDD P l=0.18u w=1.35u 
MM7 VDD B2 7 VDD P l=0.185493u w=1.42u 
MM6 VDD 6 Z VDD P l=0.186094u w=1.28u 
MM4 Z 6 VSS VSS N l=0.188166u w=1.014u 
MM3 6 A1 10 VSS N l=0.18u w=1.01u 
MM2 6 B1 11 VSS N l=0.18u w=1.01u 
MM5 10 A2 VSS VSS N l=0.18u w=1.01u 
MM1 VSS B2 11 VSS N l=0.189101u w=1.101u 
.ENDS aor22d1

.SUBCKT aor22d2 Z  A1 A2 B1 B2 VDD VSS
MM12 7 A2 6 VDD P l=0.18u w=1.35u 
MM11 7 A1 6 VDD P l=0.185815u w=1.424u 
MM10 VDD B1 7 VDD P l=0.18u w=1.35u 
MM9 VDD B2 7 VDD P l=0.185493u w=1.42u 
MM8 VDD 6 Z VDD P l=0.186142u w=1.27u 
MM7 VDD 6 Z VDD P l=0.18u w=1.2u 
MM5 Z 6 VSS VSS N l=0.187569u w=1.094u 
MM4 Z 6 VSS VSS N l=0.18u w=0.94u 
MM3 6 A1 10 VSS N l=0.18u w=1.01u 
MM2 6 B1 11 VSS N l=0.18u w=1.01u 
MM6 10 A2 VSS VSS N l=0.18u w=1.01u 
MM1 VSS B2 11 VSS N l=0.189101u w=1.101u 
.ENDS aor22d2

.SUBCKT aor22d4 Z  A1 A2 B1 B2 VDD VSS
MM14 9 A2 6 VDD P l=0.18u w=1.35u 
MM13 9 A1 6 VDD P l=0.185815u w=1.424u 
MM12 VDD B1 9 VDD P l=0.18u w=1.35u 
MM11 VDD B2 9 VDD P l=0.185493u w=1.42u 
MM10 VDD 6 Z VDD P l=0.183786u w=2.06u 
MM9 VDD 6 Z VDD P l=0.18u w=1.99u 
MM8 VDD 6 Z VDD P l=0.18u w=1.99u 
MM6 Z 6 VSS VSS N l=0.184917u w=1.684u 
MM5 Z 6 VSS VSS N l=0.18u w=1.61u 
MM4 VSS 6 Z VSS N l=0.18u w=1.61u 
MM3 6 A1 10 VSS N l=0.18u w=0.94u 
MM2 6 B1 11 VSS N l=0.18u w=1.01u 
MM7 VSS A2 10 VSS N l=0.18u w=0.94u 
MM1 VSS B2 11 VSS N l=0.189101u w=1.101u 
.ENDS aor22d4

.SUBCKT aor311d1 Z  A B C1 C2 C3 VDD VSS
MM12 VDD 2 Z VDD P l=0.18u w=1.37u 
MM11 8 C3 VDD VDD P l=0.185734u w=1.444u 
MM10 8 C2 VDD VDD P l=0.18u w=1.37u 
MM9 8 C1 VDD VDD P l=0.18u w=1.37u 
MM8 8 B 13 VDD P l=0.185417u w=1.44u 
MM7 2 A 13 VDD P l=0.185417u w=1.44u 
MM6 Z 2 VSS VSS N l=0.18u w=1.15u 
MM5 11 C3 VSS VSS N l=0.18u w=0.79u 
MM4 11 C2 12 VSS N l=0.18u w=0.79u 
MM3 2 C1 12 VSS N l=0.18u w=0.79u 
MM2 2 B VSS VSS N l=0.185738u w=1.192u 
MM1 2 A VSS VSS N l=0.18612u w=1.196u 
.ENDS aor311d1

.SUBCKT aor311d2 Z  A B C1 C2 C3 VDD VSS
MM13 VDD 3 Z VDD P l=0.185417u w=1.44u 
MM12 VDD 3 Z VDD P l=0.18u w=1.37u 
MM14 8 C2 VDD VDD P l=0.18u w=1.37u 
MM11 8 C3 VDD VDD P l=0.185734u w=1.444u 
MM10 8 C1 VDD VDD P l=0.18u w=1.37u 
MM9 8 B 13 VDD P l=0.185417u w=1.44u 
MM8 3 A 13 VDD P l=0.185417u w=1.44u 
MM6 Z 3 VSS VSS N l=0.186393u w=1.22u 
MM5 Z 3 VSS VSS N l=0.18u w=1.15u 
MM7 11 C2 12 VSS N l=0.18u w=0.79u 
MM4 11 C3 VSS VSS N l=0.18u w=0.79u 
MM3 3 C1 12 VSS N l=0.18u w=0.79u 
MM2 3 B VSS VSS N l=0.185738u w=1.192u 
MM1 3 A VSS VSS N l=0.18612u w=1.196u 
.ENDS aor311d2

.SUBCKT aor311d4 Z  A B C1 C2 C3 VDD VSS
MM16 VDD 2 Z VDD P l=0.184152u w=1.994u 
MM15 VDD 2 Z VDD P l=0.18u w=1.8u 
MM14 VDD 2 Z VDD P l=0.18u w=1.92u 
MM12 8 B 13 VDD P l=0.18u w=1.04u 
MM9 8 C1 VDD VDD P l=0.18u w=1.8u 
MM11 2 A 13 VDD P l=0.18u w=1.04u 
MM13 VDD C3 8 VDD P l=0.18u w=1.8u 
MM10 8 C2 VDD VDD P l=0.183673u w=1.862u 
MM8 VSS 2 Z VSS N l=0.18u w=1.15u 
MM7 VSS 2 Z VSS N l=0.186765u w=1.224u 
MM6 VSS 2 Z VSS N l=0.186393u w=1.22u 
MM3 2 A VSS VSS N l=0.18u w=0.76u 
MM5 11 C3 VSS VSS N l=0.18u w=1.23u 
MM2 11 C2 12 VSS N l=0.18u w=1.23u 
MM4 VSS B 2 VSS N l=0.186559u w=1.116u 
MM1 12 C1 2 VSS N l=0.18u w=1.23u 
.ENDS aor311d4

.SUBCKT aor31d1 Z  A B1 B2 B3 VDD VSS
MM8 Z 4 VDD VDD P l=0.185732u w=1.612u 
MM10 VDD B2 7 VDD P l=0.186877u w=1.204u 
MM9 VDD B3 7 VDD P l=0.18u w=1.13u 
MM7 7 B1 VDD VDD P l=0.18u w=1.13u 
MM6 4 A 7 VDD P l=0.1865u w=1.2u 
MM5 10 B2 11 VSS N l=0.18u w=1.03u 
MM4 10 B3 VSS VSS N l=0.186264u w=1.092u 
MM3 VSS 4 Z VSS N l=0.18u w=0.96u 
MM2 11 B1 4 VSS N l=0.1875u w=1.104u 
MM1 VSS A 4 VSS N l=0.186322u w=1.082u 
.ENDS aor31d1

.SUBCKT aor31d2 Z  A B1 B2 B3 VDD VSS
MM11 Z 3 VDD VDD P l=0.184407u w=1.77u 
MM10 VDD 3 Z VDD P l=0.18u w=1.7u 
MM12 VDD B3 7 VDD P l=0.18u w=1.05u 
MM9 VDD B2 7 VDD P l=0.186559u w=1.116u 
MM8 VDD B1 7 VDD P l=0.18u w=1.14u 
MM7 3 A 7 VDD P l=0.186446u w=1.21u 
MM5 VSS 3 Z VSS N l=0.18661u w=1.18u 
MM4 Z 3 VSS VSS N l=0.18u w=1.11u 
MM6 10 B3 VSS VSS N l=0.186322u w=1.082u 
MM3 10 B2 11 VSS N l=0.18u w=1.02u 
MM2 11 B1 3 VSS N l=0.187569u w=1.094u 
MM1 VSS A 3 VSS N l=0.186322u w=1.082u 
.ENDS aor31d2

.SUBCKT aor31d4 Z  A B1 B2 B3 VDD VSS
MM14 Z 2 VDD VDD P l=0.183786u w=2.06u 
MM13 Z 2 VDD VDD P l=0.18u w=1.99u 
MM12 Z 2 VDD VDD P l=0.183786u w=2.06u 
MM11 VDD B3 9 VDD P l=0.18u w=1.05u 
MM10 VDD B2 9 VDD P l=0.186559u w=1.116u 
MM9 VDD B1 9 VDD P l=0.18u w=1.14u 
MM8 2 A 9 VDD P l=0.186446u w=1.21u 
MM6 VSS 2 Z VSS N l=0.184643u w=1.68u 
MM7 VSS 2 Z VSS N l=0.184643u w=1.68u 
MM5 VSS 2 Z VSS N l=0.18u w=1.61u 
MM4 VSS B3 10 VSS N l=0.186322u w=1.082u 
MM3 10 B2 11 VSS N l=0.18u w=1.02u 
MM2 11 B1 2 VSS N l=0.187569u w=1.094u 
MM1 VSS A 2 VSS N l=0.186322u w=1.082u 
.ENDS aor31d4

.SUBCKT bh01d1   I VDD VSS
MM12 24 2 I VDD P l=0.180u w=0.420u
MM13 20 2 VDD VDD P l=0.180u w=0.420u
MM10 21 2 20 VDD P l=0.180u w=0.420u
MM9 22 2 21 VDD P l=0.180u w=0.420u
MM14 23 2 22 VDD P l=0.180u w=0.420u
MM11 24 2 23 VDD P l=0.180u w=0.420u
MM8 2 I VDD VDD P l=0.180u w=0.720u
MM1 2 I VSS VSS N l=0.180u w=0.430u
MM2 17 2 I VSS N l=0.180u w=0.300u
MM7 13 2 VSS VSS N l=0.180u w=0.300u
MM6 14 2 13 VSS N l=0.180u w=0.300u
MM5 15 2 14 VSS N l=0.180u w=0.300u
MM4 16 2 15 VSS N l=0.180u w=0.300u
MM3 17 2 16 VSS N l=0.180u w=0.300u
.ENDS bh01d1

.SUBCKT bufbd1 Z  I VDD VSS
MM5 Z 2 VDD VDD P l=0.186877u w=1.204u 
MM4 Z 2 VDD VDD P l=0.18u w=1.13u 
MM3 2 I VDD VDD P l=0.1865u w=1.2u 
MM2 VSS 2 Z VSS N l=0.18u w=0.84u 
MM1 VSS I 2 VSS N l=0.18u w=0.5u 
.ENDS bufbd1

.SUBCKT bufbd3 Z  I VDD VSS
MM8 VDD 2 Z VDD P l=0.184395u w=1.884u 
MM7 VDD 2 Z VDD P l=0.18u w=1.81u 
MM6 VDD 2 Z VDD P l=0.184395u w=1.884u 
MM5 2 I VDD VDD P l=0.186115u w=1.354u 
MM4 2 I VDD VDD P l=0.18u w=1.28u 
MM3 VSS 2 Z VSS N l=0.18u w=1.29u 
MM2 VSS 2 Z VSS N l=0.18607u w=1.364u 
MM1 2 I VSS VSS N l=0.18u w=1u 
.ENDS bufbd3

.SUBCKT bufbd7 Z  I VDD VSS
MM16 Z 2 VDD VDD P l=0.184565u w=1.814u 
MM15 Z 2 VDD VDD P l=0.184803u w=1.724u 
MM14 Z 2 VDD VDD P l=0.18u w=1.74u 
MM13 Z 2 VDD VDD P l=0.184565u w=1.814u 
MM12 VDD 2 Z VDD P l=0.18u w=1.74u 
MM11 VDD 2 Z VDD P l=0.184565u w=1.814u 
MM10 Z 2 VDD VDD P l=0.18u w=1.74u 
MM8 2 I VDD VDD P l=0.184494u w=1.522u 
MM9 VDD I 2 VDD P l=0.184436u w=1.542u 
MM7 VDD I 2 VDD P l=0.184436u w=1.542u 
MM6 Z 2 VSS VSS N l=0.186193u w=1.492u 
MM5 VSS 2 Z VSS N l=0.18u w=1.41u 
MM4 Z 2 VSS VSS N l=0.186193u w=1.492u 
MM3 Z 2 VSS VSS N l=0.18u w=0.99u 
MM2 VSS I 2 VSS N l=0.18u w=0.8u 
MM1 2 I VSS VSS N l=0.18u w=0.8u 
.ENDS bufbd7

.SUBCKT bufbda Z  I VDD VSS
MM19 VDD 2 Z VDD P l=0.184132u w=2.004u 
MM18 VDD 2 Z VDD P l=0.18u w=1.93u 
MM20 Z 2 VDD VDD P l=0.184132u w=2.004u 
MM17 Z 2 VDD VDD P l=0.18u w=1.93u 
MM16 Z 2 VDD VDD P l=0.183434u w=1.992u 
MM15 Z 2 VDD VDD P l=0.18u w=1.93u 
MM14 VDD 2 Z VDD P l=0.18u w=1.93u 
MM11 VDD 2 Z VDD P l=0.184304u w=1.924u 
MM13 Z 2 VDD VDD P l=0.184539u w=1.824u 
MM12 Z 2 VDD VDD P l=0.18u w=1.75u 
MM9 2 I VDD VDD P l=0.184524u w=1.512u 
MM10 2 I VDD VDD P l=0.184407u w=1.552u 
MM8 2 I VDD VDD P l=0.18u w=1.49u 
MM7 VSS 2 Z VSS N l=0.188404u w=1.742u 
MM6 VSS 2 Z VSS N l=0.185731u w=1.696u 
MM5 Z 2 VSS VSS N l=0.18669u w=1.713u 
MM2 VSS I 2 VSS N l=0.18u w=0.8u 
MM1 2 I VSS VSS N l=0.18u w=0.8u 
MM4 VSS 2 Z VSS N l=0.188404u w=1.742u 
MM3 Z 2 VSS VSS N l=0.185461u w=1.692u 
.ENDS bufbda

.SUBCKT buffd1 Z  I VDD VSS
MM4 VDD 2 Z VDD P l=0.184615u w=1.482u 
MM3 VDD I 2 VDD P l=0.18u w=0.57u 
MM2 Z 2 VSS VSS N l=0.186444u w=1.136u 
MM1 2 I VSS VSS N l=0.18u w=0.51u 
.ENDS buffd1

.SUBCKT buffd3 Z  I VDD VSS
MM6 VDD 2 Z VDD P l=0.184012u w=2.064u 
MM5 VDD 2 Z VDD P l=0.18u w=1.99u 
MM4 VDD I 2 VDD P l=0.18u w=1u 
MM3 VSS 2 Z VSS N l=0.18558u w=1.484u 
MM2 VSS 2 Z VSS N l=0.18u w=1.41u 
MM1 2 I VSS VSS N l=0.18u w=0.8u 
.ENDS buffd3

.SUBCKT buffd7 Z  I VDD VSS
MM12 VDD 2 Z VDD P l=0.18335u w=2.042u 
MM11 VDD 2 Z VDD P l=0.18335u w=2.042u 
MM10 Z 2 VDD VDD P l=0.18335u w=2.042u 
MM13 VDD 2 Z VDD P l=0.18335u w=2.042u 
MM9 VDD 2 Z VDD P l=0.18335u w=2.042u 
MM8 2 I VDD VDD P l=0.186u w=1.3u 
MM7 2 I VDD VDD P l=0.18u w=1.23u 
MM6 Z 2 VSS VSS N l=0.18u w=1.61u 
MM5 Z 2 VSS VSS N l=0.18u w=1.61u 
MM4 VSS 2 Z VSS N l=0.18u w=1.61u 
MM3 VSS 2 Z VSS N l=0.18u w=1.61u 
MM2 VSS I 2 VSS N l=0.18u w=0.88u 
MM1 2 I VSS VSS N l=0.18u w=0.88u 
.ENDS buffd7

.SUBCKT buffda Z  I VDD VSS
MM19 Z 2 VDD VDD P l=0.18335u w=2.042u 
MM17 VDD 2 Z VDD P l=0.18u w=1.98u 
MM16 VDD 2 Z VDD P l=0.184031u w=2.054u 
MM15 VDD 2 Z VDD P l=0.18u w=1.98u 
MM14 Z 2 VDD VDD P l=0.18335u w=2.042u 
MM18 Z 2 VDD VDD P l=0.184031u w=2.054u 
MM13 Z 2 VDD VDD P l=0.18u w=1.98u 
MM12 VDD I 2 VDD P l=0.186u w=1.3u 
MM11 VDD I 2 VDD P l=0.185294u w=1.292u 
MM10 2 I VDD VDD P l=0.18u w=1.23u 
MM9 VSS 2 Z VSS N l=0.18u w=1.61u 
MM8 VSS 2 Z VSS N l=0.18u w=1.61u 
MM7 VSS 2 Z VSS N l=0.18u w=1.61u 
MM6 VSS 2 Z VSS N l=0.18u w=1.61u 
MM5 VSS 2 Z VSS N l=0.18u w=1.61u 
MM4 Z 2 VSS VSS N l=0.18u w=1.61u 
MM3 2 I VSS VSS N l=0.18u w=0.88u 
MM2 VSS I 2 VSS N l=0.18u w=0.88u 
MM1 VSS I 2 VSS N l=0.18u w=0.88u 
.ENDS buffda

.SUBCKT buftd1 Z  EN I VDD VSS
MM9 6 EN 4 VDD P l=0.18u w=1.05u 
MM10 VDD 2 4 VDD P l=0.18u w=1.05u 
MM8 2 EN VDD VDD P l=0.18u w=0.65u 
MM7 Z 4 VDD VDD P l=0.18u w=1.56u 
MM6 4 I VDD VDD P l=0.184217u w=1.622u 
MM5 4 2 6 VSS N l=0.189854u w=1.163u 
MM4 VSS EN 2 VSS N l=0.18u w=0.52u 
MM3 VSS EN 6 VSS N l=0.18u w=1.06u 
MM2 VSS 6 Z VSS N l=0.18u w=1.03u 
MM1 VSS I 6 VSS N l=0.186264u w=1.092u 
.ENDS buftd1

.SUBCKT buftd2 Z  EN I VDD VSS
MM12 Z 2 VDD VDD P l=0.184217u w=1.622u 
MM11 Z 2 VDD VDD P l=0.18u w=1.56u 
MM10 2 I VDD VDD P l=0.184217u w=1.622u 
MM8 6 EN 2 VDD P l=0.18u w=1.05u 
MM9 VDD 4 2 VDD P l=0.18u w=1.05u 
MM7 4 EN VDD VDD P l=0.18u w=0.65u 
MM6 Z 6 VSS VSS N l=0.186096u w=1.122u 
MM5 VSS 6 Z VSS N l=0.18u w=1.06u 
MM4 VSS I 6 VSS N l=0.186096u w=1.122u 
MM3 2 4 6 VSS N l=0.189854u w=1.163u 
MM2 VSS EN 6 VSS N l=0.187302u w=1.134u 
MM1 VSS EN 4 VSS N l=0.18u w=0.52u 
.ENDS buftd2

.SUBCKT buftd4 Z  EN I VDD VSS
MM14 VDD I 3 VDD P l=0.184785u w=1.63u 
MM13 Z 3 VDD VDD P l=0.184152u w=1.994u 
MM12 Z 3 VDD VDD P l=0.18u w=1.92u 
MM11 Z 3 VDD VDD P l=0.18u w=1.92u 
MM10 VDD 4 3 VDD P l=0.18u w=1.05u 
MM9 6 EN 3 VDD P l=0.186559u w=1.116u 
MM8 4 EN VDD VDD P l=0.18u w=0.65u 
MM7 Z 6 VSS VSS N l=0.186026u w=1.374u 
MM6 Z 6 VSS VSS N l=0.18u w=1.3u 
MM5 Z 6 VSS VSS N l=0.18u w=1.3u 
MM4 VSS I 6 VSS N l=0.186207u w=1.102u 
MM3 3 4 6 VSS N l=0.187302u w=1.134u 
MM2 VSS EN 6 VSS N l=0.18u w=1.06u 
MM1 VSS EN 4 VSS N l=0.18u w=0.52u 
.ENDS buftd4

.SUBCKT buftd7 Z  EN I VDD VSS
MM18 Z 2 VDD VDD P l=0.184152u w=1.994u 
MM17 Z 2 VDD VDD P l=0.18u w=1.92u 
MM16 Z 2 VDD VDD P l=0.18u w=1.92u 
MM15 Z 2 VDD VDD P l=0.184152u w=1.994u 
MM14 Z 2 VDD VDD P l=0.18u w=1.92u 
MM13 VDD I 2 VDD P l=0.184432u w=1.76u 
MM12 VDD 4 2 VDD P l=0.18u w=1.05u 
MM11 6 EN 2 VDD P l=0.186559u w=1.116u 
MM10 4 EN VDD VDD P l=0.18u w=0.65u 
MM9 Z 6 VSS VSS N l=0.186026u w=1.374u 
MM7 VSS 6 Z VSS N l=0.18u w=1.3u 
MM8 VSS 6 Z VSS N l=0.186026u w=1.374u 
MM6 Z 6 VSS VSS N l=0.18u w=1.3u 
MM5 VSS 6 Z VSS N l=0.18u w=1.3u 
MM4 VSS I 6 VSS N l=0.185922u w=1.236u 
MM3 2 4 6 VSS N l=0.187302u w=1.134u 
MM2 VSS EN 6 VSS N l=0.18u w=1.06u 
MM1 VSS EN 4 VSS N l=0.18u w=0.52u 
.ENDS buftd7

.SUBCKT buftda Z  EN I VDD VSS
MM22 Z 2 VDD VDD P l=0.184152u w=1.994u 
MM21 Z 2 VDD VDD P l=0.18u w=1.92u 
MM20 Z 2 VDD VDD P l=0.18u w=1.92u 
MM19 Z 2 VDD VDD P l=0.184152u w=1.994u 
MM18 Z 2 VDD VDD P l=0.18u w=1.92u 
MM17 VDD 2 Z VDD P l=0.184152u w=1.994u 
MM16 Z 2 VDD VDD P l=0.18u w=1.92u 
MM15 VDD I 2 VDD P l=0.184432u w=1.76u 
MM14 VDD 4 2 VDD P l=0.18u w=1.05u 
MM13 6 EN 2 VDD P l=0.186559u w=1.116u 
MM12 4 EN VDD VDD P l=0.18u w=0.65u 
MM11 Z 6 VSS VSS N l=0.185398u w=1.534u 
MM8 VSS 6 Z VSS N l=0.18u w=1.46u 
MM10 VSS 6 Z VSS N l=0.185398u w=1.534u 
MM7 Z 6 VSS VSS N l=0.18u w=1.46u 
MM9 VSS 6 Z VSS N l=0.185398u w=1.534u 
MM6 VSS 6 Z VSS N l=0.18u w=1.46u 
MM5 Z 6 VSS VSS N l=0.18u w=1.46u 
MM4 VSS I 6 VSS N l=0.185552u w=1.232u 
MM3 2 4 6 VSS N l=0.187302u w=1.134u 
MM2 VSS EN 6 VSS N l=0.18u w=1.06u 
MM1 VSS EN 4 VSS N l=0.18u w=0.52u 
.ENDS buftda

.SUBCKT cg01d0 CO  A B CI VDD VSS
MM12 5 CI 8 VDD P l=0.18u w=1.2u 
MM11 VDD B 8 VDD P l=0.18u w=1.2u 
MM10 11 B VDD VDD P l=0.18u w=1.2u 
MM9 11 A 5 VDD P l=0.18u w=1.2u 
MM8 VDD A 8 VDD P l=0.18u w=1.2u 
MM7 VDD 5 CO VDD P l=0.18u w=0.75u 
MM6 5 CI 9 VSS N l=0.18u w=0.6u 
MM5 VSS B 9 VSS N l=0.18u w=0.6u 
MM4 VSS B 10 VSS N l=0.18u w=0.6u 
MM3 5 A 10 VSS N l=0.18u w=0.6u 
MM2 9 A VSS VSS N l=0.18u w=0.6u 
MM1 VSS 5 CO VSS N l=0.18u w=0.54u 
.ENDS cg01d0

.SUBCKT cg01d1 CO  A B CI VDD VSS
MM12 5 CI 8 VDD P l=0.18u w=1.11u 
MM11 VDD B 8 VDD P l=0.18u w=1.11u 
MM9 VDD A 8 VDD P l=0.18u w=1.11u 
MM10 11 B VDD VDD P l=0.18u w=1.11u 
MM8 11 A 5 VDD P l=0.18u w=1.11u 
MM7 VDD 5 CO VDD P l=0.18u w=1.5u 
MM6 9 CI 5 VSS N l=0.18u w=0.55u 
MM5 9 B VSS VSS N l=0.18u w=0.55u 
MM4 VSS B 10 VSS N l=0.18u w=0.55u 
MM3 10 A 5 VSS N l=0.18u w=0.55u 
MM2 VSS A 9 VSS N l=0.18u w=0.55u 
MM1 CO 5 VSS VSS N l=0.18u w=0.99u 
.ENDS cg01d1

.SUBCKT cg01d2 CO  A B CI VDD VSS
MM12 VDD A 8 VDD P l=0.18u w=1.1u 
MM13 11 B VDD VDD P l=0.18u w=1.1u 
MM11 11 A 4 VDD P l=0.18u w=1.1u 
MM10 VDD 4 CO VDD P l=0.184968u w=1.57u 
MM9 VDD 4 CO VDD P l=0.18u w=1.5u 
MM8 4 CI 8 VDD P l=0.18u w=1.1u 
MM14 VDD B 8 VDD P l=0.18u w=1.1u 
MM6 VSS B 10 VSS N l=0.18u w=0.74u 
MM5 10 A 4 VSS N l=0.18u w=0.74u 
MM4 VSS A 9 VSS N l=0.18u w=0.58u 
MM3 CO 4 VSS VSS N l=0.187569u w=1.094u 
MM2 CO 4 VSS VSS N l=0.18u w=1.02u 
MM7 9 B VSS VSS N l=0.18u w=0.58u 
MM1 9 CI 4 VSS N l=0.18u w=0.74u 
.ENDS cg01d2

.SUBCKT clk2d2 C CN  CLK VDD VSS
MM26 VDD C 9 VDD P l=0.18u w=0.57u 
MM25 VDD 3 11 VDD P l=0.18u w=0.57u 
MM24 C 4 VDD VDD P l=0.18u w=1.64u 
MM23 VDD 4 C VDD P l=0.18u w=1.64u 
MM22 VDD CN 10 VDD P l=0.18u w=0.57u 
MM21 VDD 6 12 VDD P l=0.18u w=0.6u 
MM20 CN 7 VDD VDD P l=0.184216u w=1.964u 
MM19 CN 7 VDD VDD P l=0.18u w=1.89u 
MM18 VDD 6 3 VDD P l=0.18u w=0.75u 
MM17 4 3 VDD VDD P l=0.18u w=1.07u 
MM16 7 6 VDD VDD P l=0.18u w=1.11u 
MM15 VDD CLK 6 VDD P l=0.18u w=1.11u 
MM13 VSS CLK 6 VSS N l=0.18u w=0.8u 
MM12 14 6 7 VSS N l=0.18u w=1.06u 
MM14 VSS 9 14 VSS N l=0.18u w=1.06u 
MM11 VSS 11 C VSS N l=0.18u w=0.8u 
MM10 VSS 11 C VSS N l=0.18u w=0.8u 
MM9 9 C VSS VSS N l=0.18u w=0.82u 
MM8 VSS 3 11 VSS N l=0.18u w=0.48u 
MM7 CN 12 VSS VSS N l=0.188336u w=1.166u 
MM6 CN 12 VSS VSS N l=0.18u w=1.08u 
MM5 VSS CN 10 VSS N l=0.18u w=0.48u 
MM4 VSS 6 12 VSS N l=0.18u w=0.44u 
MM2 VSS 6 3 VSS N l=0.18u w=0.57u 
MM1 4 3 15 VSS N l=0.18u w=1.03u 
MM3 VSS 10 15 VSS N l=0.18u w=1.03u 
.ENDS clk2d2

.SUBCKT cload1   I VDD VSS
MM2 VDD I VDD VDD P l=0.18u w=1.43u 
MM1 VSS I VSS VSS N l=0.18u w=0.96u 
.ENDS cload1

.SUBCKT decfq1 Q  CDN CPN D ENN VDD VSS
MM38 VDD 2 8 VDD P l=0.18u w=0.59u 
MM37 VDD CPN 2 VDD P l=0.18u w=0.59u 
MM35 VDD D 18 VDD P l=0.18u w=0.48u 
MM34 18 6 20 VDD P l=0.18u w=0.53u 
MM36 VDD 4 19 VDD P l=0.18u w=0.48u 
MM33 19 7 20 VDD P l=0.18u w=0.53u 
MM32 VDD 7 6 VDD P l=0.18u w=0.53u 
MM24 9 12 VDD VDD P l=0.18u w=0.72u 
MM21 9 8 11 VDD P l=0.18u w=0.53u 
MM31 12 2 20 VDD P l=0.18u w=0.52u 
MM30 4 2 11 VDD P l=0.18u w=0.53u 
MM27 4 10 VDD VDD P l=0.18u w=0.48u 
MM29 12 8 17 VDD P l=0.18u w=0.52u 
MM28 VDD 9 17 VDD P l=0.18u w=0.53u 
MM26 VDD 10 Q VDD P l=0.18u w=1.51u 
MM25 VDD 11 10 VDD P l=0.18u w=0.98u 
MM23 VDD CDN 10 VDD P l=0.18u w=0.98u 
MM22 VDD CDN 17 VDD P l=0.18u w=0.52u 
MM20 VDD ENN 7 VDD P l=0.18u w=0.81u 
MM17 4 8 11 VSS N l=0.18u w=0.48u 
MM14 4 10 VSS VSS N l=0.18u w=0.48u 
MM18 9 2 11 VSS N l=0.18u w=0.48u 
MM19 12 2 17 VSS N l=0.18u w=0.48u 
MM16 12 8 20 VSS N l=0.18u w=0.48u 
MM13 VSS 12 9 VSS N l=0.18u w=0.61u 
MM12 21 CDN 17 VSS N l=0.18u w=0.53u 
MM15 VSS 9 21 VSS N l=0.18u w=0.53u 
MM11 VSS 2 8 VSS N l=0.18u w=0.48u 
MM10 VSS CPN 2 VSS N l=0.18u w=0.47u 
MM7 19 6 20 VSS N l=0.18u w=0.5u 
MM5 20 7 18 VSS N l=0.18u w=0.5u 
MM9 19 4 VSS VSS N l=0.18u w=0.5u 
MM6 VSS 7 6 VSS N l=0.18u w=0.44u 
MM8 VSS D 18 VSS N l=0.18u w=0.5u 
MM4 VSS ENN 7 VSS N l=0.18u w=0.48u 
MM3 Q 10 VSS VSS N l=0.18u w=0.99u 
MM2 10 11 22 VSS N l=0.18u w=0.99u 
MM1 22 CDN VSS VSS N l=0.18u w=0.99u 
.ENDS decfq1

.SUBCKT decfq2 Q  CDN CPN D ENN VDD VSS
MM40 VDD 2 8 VDD P l=0.18u w=0.59u 
MM39 VDD CPN 2 VDD P l=0.18u w=0.59u 
MM37 VDD D 18 VDD P l=0.18u w=0.48u 
MM36 18 6 20 VDD P l=0.18u w=0.53u 
MM38 VDD 4 19 VDD P l=0.18u w=0.48u 
MM35 19 7 20 VDD P l=0.18u w=0.53u 
MM34 VDD 7 6 VDD P l=0.18u w=0.53u 
MM25 9 12 VDD VDD P l=0.18u w=0.72u 
MM22 9 8 11 VDD P l=0.18u w=0.53u 
MM33 12 2 20 VDD P l=0.18u w=0.52u 
MM32 4 2 11 VDD P l=0.18u w=0.53u 
MM29 4 10 VDD VDD P l=0.18u w=0.48u 
MM31 12 8 17 VDD P l=0.18u w=0.52u 
MM30 VDD 9 17 VDD P l=0.18u w=0.53u 
MM28 VDD 10 Q VDD P l=0.184379u w=1.562u 
MM27 VDD 10 Q VDD P l=0.184674u w=1.566u 
MM26 VDD 11 10 VDD P l=0.18u w=0.98u 
MM24 VDD CDN 10 VDD P l=0.18u w=0.98u 
MM23 VDD CDN 17 VDD P l=0.18u w=0.52u 
MM21 VDD ENN 7 VDD P l=0.18u w=0.81u 
MM18 4 8 11 VSS N l=0.18u w=0.48u 
MM15 4 10 VSS VSS N l=0.18u w=0.48u 
MM19 9 2 11 VSS N l=0.18u w=0.48u 
MM20 12 2 17 VSS N l=0.18u w=0.48u 
MM17 12 8 20 VSS N l=0.18u w=0.48u 
MM14 VSS 12 9 VSS N l=0.18u w=0.61u 
MM13 21 CDN 17 VSS N l=0.18u w=0.53u 
MM16 VSS 9 21 VSS N l=0.18u w=0.53u 
MM12 VSS 10 Q VSS N l=0.186502u w=1.052u 
MM11 Q 10 VSS VSS N l=0.186502u w=1.052u 
MM10 10 11 22 VSS N l=0.18u w=0.99u 
MM9 22 CDN VSS VSS N l=0.18u w=0.99u 
MM8 VSS 2 8 VSS N l=0.18u w=0.48u 
MM7 VSS CPN 2 VSS N l=0.18u w=0.47u 
MM4 19 6 20 VSS N l=0.18u w=0.5u 
MM2 20 7 18 VSS N l=0.18u w=0.5u 
MM6 19 4 VSS VSS N l=0.18u w=0.5u 
MM3 VSS 7 6 VSS N l=0.18u w=0.44u 
MM5 VSS D 18 VSS N l=0.18u w=0.5u 
MM1 VSS ENN 7 VSS N l=0.18u w=0.48u 
.ENDS decfq2

.SUBCKT decrq1 Q  CDN CP D ENN VDD VSS
MM37 VDD 3 12 VDD P l=0.18u w=0.49u 
MM38 3 CDN VDD VDD P l=0.18u w=1.05u 
MM36 3 4 VDD VDD P l=0.18u w=1.05u 
MM35 Q 3 VDD VDD P l=0.18u w=1.5u 
MM33 6 5 4 VDD P l=0.18u w=0.6u 
MM30 VDD 7 6 VDD P l=0.18u w=0.82u 
MM34 VDD CDN 15 VDD P l=0.18u w=0.6u 
MM32 15 5 7 VDD P l=0.18u w=0.6u 
MM31 VDD 6 15 VDD P l=0.18u w=0.6u 
MM29 12 8 4 VDD P l=0.18u w=0.6u 
MM28 20 8 7 VDD P l=0.18u w=0.6u 
MM27 8 5 VDD VDD P l=0.18u w=0.68u 
MM25 VDD CP 5 VDD P l=0.18u w=0.68u 
MM24 18 11 20 VDD P l=0.18u w=0.6u 
MM22 20 13 19 VDD P l=0.18u w=0.6u 
MM26 18 D VDD VDD P l=0.18u w=0.52u 
MM23 VDD 12 19 VDD P l=0.18u w=0.43u 
MM21 VDD ENN 13 VDD P l=0.18u w=0.93u 
MM20 11 13 VDD VDD P l=0.18u w=0.6u 
MM19 21 CDN 15 VSS N l=0.18u w=0.6u 
MM11 7 8 15 VSS N l=0.18u w=0.44u 
MM17 VSS 5 8 VSS N l=0.18u w=0.52u 
MM16 20 5 7 VSS N l=0.18u w=0.44u 
MM15 21 6 VSS VSS N l=0.18u w=0.6u 
MM18 12 5 4 VSS N l=0.18u w=0.44u 
MM14 VSS 3 12 VSS N l=0.18u w=0.44u 
MM13 VSS 7 6 VSS N l=0.18u w=0.7u 
MM12 4 8 6 VSS N l=0.18u w=0.44u 
MM10 22 CDN VSS VSS N l=0.18u w=1.05u 
MM9 22 4 3 VSS N l=0.18u w=1.05u 
MM8 Q 3 VSS VSS N l=0.18u w=1u 
MM7 VSS 13 11 VSS N l=0.18u w=0.43u 
MM6 20 13 18 VSS N l=0.18u w=0.42u 
MM5 VSS D 18 VSS N l=0.18u w=0.42u 
MM4 VSS CP 5 VSS N l=0.18u w=0.53u 
MM3 19 11 20 VSS N l=0.18u w=0.44u 
MM2 19 12 VSS VSS N l=0.18u w=0.44u 
MM1 VSS ENN 13 VSS N l=0.18u w=0.43u 
.ENDS decrq1

.SUBCKT decrq2 Q  CDN CP D ENN VDD VSS
MM38 2 4 8 VDD P l=0.18u w=0.6u 
MM36 VDD 5 2 VDD P l=0.18u w=0.82u 
MM40 VDD 2 15 VDD P l=0.18u w=0.6u 
MM39 VDD CDN 15 VDD P l=0.18u w=0.6u 
MM37 15 4 5 VDD P l=0.18u w=0.6u 
MM35 12 6 8 VDD P l=0.18u w=0.6u 
MM34 20 6 5 VDD P l=0.18u w=0.6u 
MM32 VDD 7 12 VDD P l=0.18u w=0.49u 
MM33 7 CDN VDD VDD P l=0.18u w=1.05u 
MM31 7 8 VDD VDD P l=0.18u w=1.05u 
MM30 Q 7 VDD VDD P l=0.1852u w=1.5u 
MM29 Q 7 VDD VDD P l=0.1852u w=1.5u 
MM27 VDD CP 4 VDD P l=0.18u w=0.68u 
MM26 18 11 20 VDD P l=0.18u w=0.6u 
MM24 20 13 19 VDD P l=0.18u w=0.6u 
MM28 18 D VDD VDD P l=0.18u w=0.52u 
MM25 VDD 12 19 VDD P l=0.18u w=0.43u 
MM23 VDD ENN 13 VDD P l=0.18u w=0.93u 
MM22 11 13 VDD VDD P l=0.18u w=0.6u 
MM21 6 4 VDD VDD P l=0.18u w=0.68u 
MM19 21 CDN 15 VSS N l=0.18u w=0.6u 
MM12 15 6 5 VSS N l=0.18u w=0.44u 
MM20 21 2 VSS VSS N l=0.18u w=0.6u 
MM17 VSS 4 6 VSS N l=0.18u w=0.52u 
MM16 20 4 5 VSS N l=0.18u w=0.44u 
MM18 12 4 8 VSS N l=0.18u w=0.44u 
MM15 VSS 7 12 VSS N l=0.18u w=0.44u 
MM14 VSS 5 2 VSS N l=0.18u w=0.7u 
MM13 8 6 2 VSS N l=0.18u w=0.44u 
MM11 22 CDN VSS VSS N l=0.18u w=1.05u 
MM10 22 8 7 VSS N l=0.18u w=1.05u 
MM9 Q 7 VSS VSS N l=0.18u w=1u 
MM8 VSS 7 Q VSS N l=0.18u w=1u 
MM7 VSS 13 11 VSS N l=0.18u w=0.43u 
MM6 20 13 18 VSS N l=0.18u w=0.42u 
MM5 VSS D 18 VSS N l=0.18u w=0.42u 
MM4 VSS CP 4 VSS N l=0.18u w=0.53u 
MM3 19 11 20 VSS N l=0.18u w=0.44u 
MM2 19 12 VSS VSS N l=0.18u w=0.44u 
MM1 VSS ENN 13 VSS N l=0.18u w=0.43u 
.ENDS decrq2

.SUBCKT denrq1 Q  CP D ENN VDD VSS
MM34 5 2 19 VDD P l=0.18u w=0.48u 
MM33 9 2 12 VDD P l=0.18u w=0.48u 
MM28 9 6 VDD VDD P l=0.18u w=0.48u 
MM32 12 3 4 VDD P l=0.18u w=0.48u 
MM31 5 3 15 VDD P l=0.18u w=0.48u 
MM30 VDD 4 15 VDD P l=0.18u w=0.48u 
MM29 VDD 5 4 VDD P l=0.18u w=0.51u 
MM27 VDD 3 2 VDD P l=0.18u w=0.51u 
MM26 VDD CP 3 VDD P l=0.18u w=0.51u 
MM25 19 8 17 VDD P l=0.18u w=0.48u 
MM23 VDD D 17 VDD P l=0.18u w=0.48u 
MM24 18 9 VDD VDD P l=0.18u w=0.48u 
MM22 18 11 19 VDD P l=0.18u w=0.48u 
MM21 VDD 11 8 VDD P l=0.18u w=0.48u 
MM20 VDD 12 6 VDD P l=0.189502u w=1.105u 
MM19 Q 6 VDD VDD P l=0.184554u w=1.502u 
MM18 VDD ENN 11 VDD P l=0.18u w=0.65u 
MM17 5 2 15 VSS N l=0.18u w=0.66u 
MM15 5 3 19 VSS N l=0.18u w=0.66u 
MM16 4 2 12 VSS N l=0.18u w=0.66u 
MM14 9 3 12 VSS N l=0.18u w=0.66u 
MM13 15 4 VSS VSS N l=0.18u w=0.66u 
MM12 4 5 VSS VSS N l=0.18u w=0.66u 
MM11 9 6 VSS VSS N l=0.18u w=0.66u 
MM10 VSS 3 2 VSS N l=0.18u w=0.48u 
MM9 VSS CP 3 VSS N l=0.18u w=0.48u 
MM8 18 8 19 VSS N l=0.18u w=0.66u 
MM7 18 9 VSS VSS N l=0.18u w=0.66u 
MM5 VSS 11 8 VSS N l=0.18u w=0.48u 
MM4 19 11 17 VSS N l=0.18u w=0.66u 
MM6 VSS D 17 VSS N l=0.18u w=0.66u 
MM3 VSS ENN 11 VSS N l=0.18u w=0.45u 
MM2 6 12 VSS VSS N l=0.18729u w=1.07u 
MM1 Q 6 VSS VSS N l=0.186826u w=1.002u 
.ENDS denrq1

.SUBCKT denrq2 Q  CP D ENN VDD VSS
MM36 5 2 19 VDD P l=0.18u w=0.48u 
MM35 10 2 7 VDD P l=0.18u w=0.48u 
MM30 10 6 VDD VDD P l=0.18u w=0.48u 
MM34 7 3 4 VDD P l=0.18u w=0.48u 
MM33 5 3 16 VDD P l=0.18u w=0.48u 
MM32 VDD 4 16 VDD P l=0.18u w=0.48u 
MM31 VDD 5 4 VDD P l=0.18u w=0.51u 
MM29 VDD 7 6 VDD P l=0.189502u w=1.105u 
MM28 Q 6 VDD VDD P l=0.184554u w=1.502u 
MM27 Q 6 VDD VDD P l=0.184554u w=1.502u 
MM26 VDD 3 2 VDD P l=0.18u w=0.51u 
MM25 VDD CP 3 VDD P l=0.18u w=0.51u 
MM24 19 9 17 VDD P l=0.18u w=0.48u 
MM22 VDD D 17 VDD P l=0.18u w=0.48u 
MM23 18 10 VDD VDD P l=0.18u w=0.48u 
MM21 18 12 19 VDD P l=0.18u w=0.48u 
MM20 VDD 12 9 VDD P l=0.18u w=0.48u 
MM19 VDD ENN 12 VDD P l=0.18u w=0.65u 
MM18 5 2 16 VSS N l=0.18u w=0.66u 
MM16 5 3 19 VSS N l=0.18u w=0.66u 
MM17 4 2 7 VSS N l=0.18u w=0.66u 
MM15 10 3 7 VSS N l=0.18u w=0.66u 
MM14 16 4 VSS VSS N l=0.18u w=0.66u 
MM13 4 5 VSS VSS N l=0.18u w=0.66u 
MM12 10 6 VSS VSS N l=0.18u w=0.66u 
MM11 6 7 VSS VSS N l=0.18729u w=1.07u 
MM10 VSS 6 Q VSS N l=0.187276u w=1.006u 
MM9 Q 6 VSS VSS N l=0.186826u w=1.002u 
MM8 VSS 3 2 VSS N l=0.18u w=0.48u 
MM7 VSS CP 3 VSS N l=0.18u w=0.48u 
MM6 18 9 19 VSS N l=0.18u w=0.66u 
MM5 18 10 VSS VSS N l=0.18u w=0.66u 
MM3 VSS 12 9 VSS N l=0.18u w=0.48u 
MM2 19 12 17 VSS N l=0.18u w=0.66u 
MM4 VSS D 17 VSS N l=0.18u w=0.66u 
MM1 VSS ENN 12 VSS N l=0.18u w=0.45u 
.ENDS denrq2

.SUBCKT depfq1 Q  CPN D ENN SDN VDD VSS
MM37 20 3 8 VDD P l=0.18u w=0.55u 
MM36 VDD SDN 2 VDD P l=0.18u w=0.75u 
MM38 VDD 2 17 VDD P l=0.18u w=0.55u 
MM35 17 5 8 VDD P l=0.18u w=0.55u 
MM34 7 6 VDD VDD P l=0.186501u w=1.126u 
MM33 Q 7 VDD VDD P l=0.18u w=1.13u 
MM32 VDD 7 9 VDD P l=0.18u w=0.64u 
MM31 VDD SDN 9 VDD P l=0.18u w=0.64u 
MM29 2 8 VDD VDD P l=0.18u w=0.42u 
MM28 2 5 6 VDD P l=0.18u w=0.6u 
MM30 9 3 6 VDD P l=0.18u w=0.6u 
MM26 19 10 20 VDD P l=0.18u w=0.48u 
MM25 19 D VDD VDD P l=0.18u w=0.48u 
MM24 VDD CPN 3 VDD P l=0.18u w=0.51u 
MM27 VDD 9 18 VDD P l=0.18u w=0.48u 
MM23 20 13 18 VDD P l=0.18u w=0.48u 
MM22 10 13 VDD VDD P l=0.18u w=0.48u 
MM21 VDD 3 5 VDD P l=0.18u w=0.52u 
MM20 VDD ENN 13 VDD P l=0.18u w=0.7u 
MM19 VSS 2 17 VSS N l=0.18u w=0.48u 
MM17 17 3 8 VSS N l=0.18u w=0.66u 
MM16 9 7 21 VSS N l=0.18u w=0.66u 
MM14 21 SDN VSS VSS N l=0.18u w=0.66u 
MM18 6 3 2 VSS N l=0.18u w=0.44u 
MM13 9 5 6 VSS N l=0.18u w=0.66u 
MM12 22 8 2 VSS N l=0.18u w=0.66u 
MM15 VSS SDN 22 VSS N l=0.18u w=0.66u 
MM11 8 5 20 VSS N l=0.18u w=0.66u 
MM10 VSS 3 5 VSS N l=0.18u w=0.52u 
MM9 7 6 VSS VSS N l=0.18u w=0.75u 
MM8 Q 7 VSS VSS N l=0.18u w=0.75u 
MM7 VSS 13 10 VSS N l=0.18u w=0.44u 
MM5 18 9 VSS VSS N l=0.18u w=0.45u 
MM4 18 10 20 VSS N l=0.18u w=0.44u 
MM6 20 13 19 VSS N l=0.18u w=0.44u 
MM3 VSS D 19 VSS N l=0.18u w=0.44u 
MM2 3 CPN VSS VSS N l=0.18u w=0.47u 
MM1 VSS ENN 13 VSS N l=0.18u w=0.48u 
.ENDS depfq1

.SUBCKT depfq2 Q  CPN D ENN SDN VDD VSS
MM40 8 2 20 VDD P l=0.18u w=0.55u 
MM39 VDD SDN IPM VDD P l=0.18u w=0.75u 
MM38 VDD IPM 17 VDD P l=0.18u w=0.55u 
MM37 17 5 8 VDD P l=0.18u w=0.55u 
MM36 7 IPS VDD VDD P l=0.186501u w=1.126u 
MM35 VDD 7 Q VDD P l=0.1865u w=1.2u 
MM34 VDD 7 Q VDD P l=0.18u w=1.13u 
MM33 9 7 VDD VDD P l=0.18u w=0.64u 
MM32 9 SDN VDD VDD P l=0.18u w=0.64u 
MM30 IPM 8 VDD VDD P l=0.18u w=0.42u 
MM29 IPM 5 IPS VDD P l=0.18u w=0.6u 
MM31 9 2 IPS VDD P l=0.18u w=0.6u 
MM27 19 10 20 VDD P l=0.18u w=0.48u 
MM26 19 D VDD VDD P l=0.18u w=0.48u 
MM25 VDD CPN 2 VDD P l=0.18u w=0.51u 
MM28 VDD 9 18 VDD P l=0.18u w=0.48u 
MM24 20 13 18 VDD P l=0.18u w=0.48u 
MM23 10 13 VDD VDD P l=0.18u w=0.48u 
MM22 VDD 2 5 VDD P l=0.18u w=0.52u 
MM21 VDD ENN 13 VDD P l=0.18u w=0.7u 
MM19 17 2 8 VSS N l=0.18u w=0.66u 
MM13 VSS IPM 17 VSS N l=0.18u w=0.48u 
MM20 IPS 2 IPM VSS N l=0.18u w=0.44u 
MM18 21 8 IPM VSS N l=0.18u w=0.66u 
MM16 VSS SDN 21 VSS N l=0.18u w=0.66u 
MM17 9 7 22 VSS N l=0.18u w=0.66u 
MM15 22 SDN VSS VSS N l=0.18u w=0.66u 
MM14 9 5 IPS VSS N l=0.18u w=0.66u 
MM12 8 5 20 VSS N l=0.18u w=0.66u 
MM11 VSS 2 5 VSS N l=0.18u w=0.52u 
MM10 VSS 13 10 VSS N l=0.18u w=0.44u 
MM8 18 9 VSS VSS N l=0.18u w=0.45u 
MM7 18 10 20 VSS N l=0.18u w=0.44u 
MM9 20 13 19 VSS N l=0.18u w=0.44u 
MM6 VSS D 19 VSS N l=0.18u w=0.44u 
MM5 2 CPN VSS VSS N l=0.18u w=0.47u 
MM4 7 IPS VSS VSS N l=0.18u w=0.79u 
MM3 VSS 7 Q VSS N l=0.18u w=0.82u 
MM2 Q 7 VSS VSS N l=0.18u w=0.82u 
MM1 VSS ENN 13 VSS N l=0.18u w=0.48u 
.ENDS depfq2

.SUBCKT deprq1 Q  CP D ENN SDN VDD VSS
MM38 5 2 19 VDD P l=0.18u w=0.48u 
MM37 5 3 16 VDD P l=0.18u w=0.48u 
MM36 VDD 4 16 VDD P l=0.18u w=0.48u 
MM35 VDD 5 4 VDD P l=0.18u w=0.57u 
MM34 VDD SDN 4 VDD P l=0.18u w=0.57u 
MM33 8 7 VDD VDD P l=0.186441u w=1.062u 
MM32 VDD 8 9 VDD P l=0.18u w=0.65u 
MM31 VDD SDN 9 VDD P l=0.18u w=0.65u 
MM29 20 10 19 VDD P l=0.18u w=0.52u 
MM28 VDD D 20 VDD P l=0.18u w=0.52u 
MM27 VDD 12 10 VDD P l=0.18u w=0.51u 
MM30 VDD 9 18 VDD P l=0.18u w=0.48u 
MM26 18 12 19 VDD P l=0.18u w=0.52u 
MM25 VDD 3 2 VDD P l=0.18u w=0.51u 
MM24 VDD CP 3 VDD P l=0.18u w=0.64u 
MM23 VDD ENN 12 VDD P l=0.18u w=0.83u 
MM22 Q 8 VDD VDD P l=0.1852u w=1.5u 
MM21 7 2 9 VDD P l=0.18u w=0.48u 
MM20 7 3 4 VDD P l=0.18u w=0.48u 
MM18 5 2 16 VSS N l=0.18u w=0.66u 
MM15 16 4 VSS VSS N l=0.18u w=0.48u 
MM17 5 3 19 VSS N l=0.18u w=0.66u 
MM16 9 3 7 VSS N l=0.18u w=0.66u 
MM13 9 8 22 VSS N l=0.18u w=0.66u 
MM19 4 2 7 VSS N l=0.18u w=0.66u 
MM14 4 5 21 VSS N l=0.18u w=0.66u 
MM12 VSS SDN 21 VSS N l=0.18u w=0.66u 
MM11 VSS SDN 22 VSS N l=0.18u w=0.66u 
MM10 18 9 VSS VSS N l=0.18u w=0.43u 
MM9 18 10 19 VSS N l=0.18u w=0.43u 
MM7 VSS 12 10 VSS N l=0.18u w=0.57u 
MM6 19 12 20 VSS N l=0.18u w=0.43u 
MM8 VSS D 20 VSS N l=0.18u w=0.43u 
MM5 VSS 3 2 VSS N l=0.18u w=0.49u 
MM4 VSS CP 3 VSS N l=0.18u w=0.49u 
MM3 VSS ENN 12 VSS N l=0.18u w=0.48u 
MM2 Q 8 VSS VSS N l=0.18u w=1u 
MM1 8 7 VSS VSS N l=0.18u w=1u 
.ENDS deprq1

.SUBCKT deprq2 Q  CP D ENN SDN VDD VSS
MM40 5 2 19 VDD P l=0.18u w=0.48u 
MM39 5 3 15 VDD P l=0.18u w=0.48u 
MM38 VDD 4 15 VDD P l=0.18u w=0.48u 
MM37 VDD 5 4 VDD P l=0.18u w=0.57u 
MM36 VDD SDN 4 VDD P l=0.18u w=0.57u 
MM35 8 7 VDD VDD P l=0.186441u w=1.062u 
MM34 10 8 VDD VDD P l=0.18u w=0.65u 
MM33 VDD SDN 10 VDD P l=0.18u w=0.65u 
MM32 VDD 3 2 VDD P l=0.18u w=0.51u 
MM31 VDD CP 3 VDD P l=0.18u w=0.64u 
MM29 20 11 19 VDD P l=0.18u w=0.52u 
MM28 VDD D 20 VDD P l=0.18u w=0.52u 
MM27 VDD 13 11 VDD P l=0.18u w=0.51u 
MM30 VDD 10 18 VDD P l=0.18u w=0.48u 
MM26 18 13 19 VDD P l=0.18u w=0.52u 
MM25 VDD ENN 13 VDD P l=0.18u w=0.83u 
MM24 Q 8 VDD VDD P l=0.185098u w=1.53u 
MM23 Q 8 VDD VDD P l=0.18u w=1.46u 
MM22 7 2 10 VDD P l=0.18u w=0.48u 
MM21 7 3 4 VDD P l=0.18u w=0.48u 
MM19 5 2 15 VSS N l=0.18u w=0.66u 
MM16 15 4 VSS VSS N l=0.18u w=0.48u 
MM18 5 3 19 VSS N l=0.18u w=0.66u 
MM17 10 3 7 VSS N l=0.18u w=0.66u 
MM14 10 8 22 VSS N l=0.18u w=0.66u 
MM20 4 2 7 VSS N l=0.18u w=0.66u 
MM15 4 5 21 VSS N l=0.18u w=0.66u 
MM13 VSS SDN 21 VSS N l=0.18u w=0.66u 
MM12 VSS SDN 22 VSS N l=0.18u w=0.66u 
MM11 Q 8 VSS VSS N l=0.187856u w=1.054u 
MM10 Q 8 VSS VSS N l=0.18u w=0.98u 
MM9 VSS 7 8 VSS N l=0.18u w=0.98u 
MM8 18 10 VSS VSS N l=0.18u w=0.43u 
MM7 18 11 19 VSS N l=0.18u w=0.43u 
MM5 VSS 13 11 VSS N l=0.18u w=0.57u 
MM4 19 13 20 VSS N l=0.18u w=0.43u 
MM6 VSS D 20 VSS N l=0.18u w=0.43u 
MM3 VSS 3 2 VSS N l=0.18u w=0.49u 
MM2 VSS CP 3 VSS N l=0.18u w=0.49u 
MM1 VSS ENN 13 VSS N l=0.18u w=0.48u 
.ENDS deprq2

.SUBCKT dfbfb1 Q QN  CDN CPN D SDN VDD VSS
MM33 10 SDN VDD VDD P l=0.18u w=0.95u 
MM29 10 6 IPS VDD P l=0.18u w=0.67u 
MM32 15 3 IPS VDD P l=0.18u w=0.73u 
MM34 15 SDN VDD VDD P l=0.187952u w=1.162u 
MM31 15 4 VDD VDD P l=0.185886u w=1.162u 
MM30 10 IPM VDD VDD P l=0.191073u w=1.165u 
MM28 VDD CDN 4 VDD P l=0.184844u w=1.412u 
MM27 VDD IPS 4 VDD P l=0.18u w=1.26u 
MM26 16 CDN VDD VDD P l=0.18u w=0.86u 
MM22 16 6 IPM VDD P l=0.18u w=0.65u 
MM25 17 3 IPM VDD P l=0.18u w=0.65u 
MM24 17 D VDD VDD P l=0.18u w=0.54u 
MM23 16 10 VDD VDD P l=0.187709u w=1.074u 
MM21 Q 4 VDD VDD P l=0.18u w=1.4u 
MM20 QN IPS VDD VDD P l=0.185306u w=1.47u 
MM19 VDD 3 6 VDD P l=0.18u w=0.68u 
MM18 VDD CPN 3 VDD P l=0.18u w=0.7u 
MM17 20 SDN 10 VSS N l=0.18u w=0.9u 
MM12 IPS 3 10 VSS N l=0.18u w=0.76u 
MM15 21 CDN 16 VSS N l=0.18u w=0.86u 
MM13 IPM 3 16 VSS N l=0.18u w=0.48u 
MM11 IPM 6 17 VSS N l=0.18u w=0.48u 
MM16 18 SDN 15 VSS N l=0.18u w=0.76u 
MM10 IPS 6 15 VSS N l=0.18u w=0.76u 
MM9 18 4 VSS VSS N l=0.18u w=0.76u 
MM8 4 IPS 19 VSS N l=0.18u w=1.07u 
MM14 VSS CDN 19 VSS N l=0.18u w=1.07u 
MM7 17 D VSS VSS N l=0.18u w=0.48u 
MM6 20 IPM VSS VSS N l=0.18u w=0.9u 
MM5 21 10 VSS VSS N l=0.18u w=0.86u 
MM4 VSS 4 Q VSS N l=0.18u w=1.06u 
MM3 VSS IPS QN VSS N l=0.186903u w=1.13u 
MM2 VSS 3 6 VSS N l=0.18u w=0.52u 
MM1 VSS CPN 3 VSS N l=0.18u w=0.52u 
.ENDS dfbfb1

.SUBCKT dfbfb2 Q QN  CDN CPN D SDN VDD VSS
MM37 10 SDN VDD VDD P l=0.18u w=0.95u 
MM35 10 4 IPS VDD P l=0.18u w=0.67u 
MM36 14 3 IPS VDD P l=0.18u w=0.73u 
MM38 14 SDN VDD VDD P l=0.187952u w=1.162u 
MM34 14 5 VDD VDD P l=0.185886u w=1.162u 
MM33 10 IPM VDD VDD P l=0.191073u w=1.165u 
MM31 QN IPS VDD VDD P l=0.18u w=1.54u 
MM30 QN IPS VDD VDD P l=0.18u w=1.54u 
MM29 VDD 5 Q VDD P l=0.18u w=1.54u 
MM28 Q 5 VDD VDD P l=0.18u w=1.54u 
MM32 VDD CDN 5 VDD P l=0.184844u w=1.412u 
MM27 VDD IPS 5 VDD P l=0.184494u w=1.522u 
MM26 16 CDN VDD VDD P l=0.18u w=0.86u 
MM22 16 4 IPM VDD P l=0.18u w=0.65u 
MM25 17 3 IPM VDD P l=0.18u w=0.65u 
MM24 17 D VDD VDD P l=0.18u w=0.54u 
MM23 16 10 VDD VDD P l=0.187709u w=1.074u 
MM21 VDD 3 4 VDD P l=0.18u w=0.68u 
MM20 VDD CPN 3 VDD P l=0.18u w=0.7u 
MM19 20 SDN 10 VSS N l=0.18u w=0.9u 
MM14 IPS 3 10 VSS N l=0.18u w=0.76u 
MM17 21 CDN 16 VSS N l=0.18u w=0.86u 
MM15 IPM 3 16 VSS N l=0.18u w=0.48u 
MM13 IPM 4 17 VSS N l=0.18u w=0.48u 
MM18 18 SDN 14 VSS N l=0.18u w=0.76u 
MM12 IPS 4 14 VSS N l=0.18u w=0.76u 
MM11 18 5 VSS VSS N l=0.18u w=0.76u 
MM10 5 IPS 19 VSS N l=0.18u w=1.07u 
MM16 VSS CDN 19 VSS N l=0.18u w=1.07u 
MM9 17 D VSS VSS N l=0.18u w=0.48u 
MM8 20 IPM VSS VSS N l=0.18u w=0.9u 
MM7 21 10 VSS VSS N l=0.18u w=0.86u 
MM6 VSS IPS QN VSS N l=0.18u w=1u 
MM5 VSS IPS QN VSS N l=0.18u w=1u 
MM4 VSS 5 Q VSS N l=0.18u w=1u 
MM3 VSS 5 Q VSS N l=0.18u w=1u 
MM2 VSS 3 4 VSS N l=0.18u w=0.52u 
MM1 VSS CPN 3 VSS N l=0.18u w=0.52u 
.ENDS dfbfb2

.SUBCKT dfbrb1 Q QN  CDN CP D SDN VDD VSS
MM34 15 2 IPS VDD P l=0.18u w=0.73u 
MM29 10 6 IPS VDD P l=0.18u w=0.67u 
MM33 15 SDN VDD VDD P l=0.187952u w=1.162u 
MM32 10 SDN VDD VDD P l=0.18u w=0.95u 
MM31 15 4 VDD VDD P l=0.185886u w=1.162u 
MM30 10 IPM VDD VDD P l=0.191073u w=1.165u 
MM28 VDD CDN 4 VDD P l=0.184844u w=1.412u 
MM27 VDD IPS 4 VDD P l=0.18u w=1.26u 
MM26 16 CDN VDD VDD P l=0.18u w=0.86u 
MM23 16 6 IPM VDD P l=0.18u w=0.65u 
MM25 17 2 IPM VDD P l=0.18u w=0.65u 
MM24 17 D VDD VDD P l=0.18u w=0.54u 
MM22 16 10 VDD VDD P l=0.187709u w=1.074u 
MM21 Q 4 VDD VDD P l=0.18u w=1.4u 
MM20 QN IPS VDD VDD P l=0.185306u w=1.47u 
MM19 VDD 6 2 VDD P l=0.18u w=0.68u 
MM18 VDD CP 6 VDD P l=0.18u w=0.7u 
MM17 IPS 2 10 VSS N l=0.18u w=0.76u 
MM15 IPS 6 15 VSS N l=0.18u w=0.76u 
MM14 20 SDN 10 VSS N l=0.18u w=0.9u 
MM13 18 SDN 15 VSS N l=0.18u w=0.76u 
MM16 IPM 2 16 VSS N l=0.18u w=0.48u 
MM12 21 CDN 16 VSS N l=0.18u w=0.86u 
MM10 18 4 VSS VSS N l=0.18u w=0.76u 
MM9 4 IPS 19 VSS N l=0.18u w=1.07u 
MM11 VSS CDN 19 VSS N l=0.18u w=1.07u 
MM7 IPM 6 17 VSS N l=0.18u w=0.48u 
MM8 17 D VSS VSS N l=0.18u w=0.48u 
MM6 20 IPM VSS VSS N l=0.18u w=0.9u 
MM5 21 10 VSS VSS N l=0.18u w=0.86u 
MM4 VSS 4 Q VSS N l=0.18u w=1.06u 
MM3 VSS IPS QN VSS N l=0.186903u w=1.13u 
MM2 VSS 6 2 VSS N l=0.18u w=0.52u 
MM1 VSS CP 6 VSS N l=0.18u w=0.52u 
.ENDS dfbrb1

.SUBCKT dfbrb2 Q QN  CDN CP D SDN VDD VSS
MM38 14 2 IPS VDD P l=0.18u w=0.73u 
MM35 10 4 IPS VDD P l=0.18u w=0.67u 
MM37 14 SDN VDD VDD P l=0.187952u w=1.162u 
MM36 10 SDN VDD VDD P l=0.18u w=0.95u 
MM34 14 5 VDD VDD P l=0.185886u w=1.162u 
MM33 10 IPM VDD VDD P l=0.191073u w=1.165u 
MM31 QN IPS VDD VDD P l=0.18u w=1.54u 
MM30 QN IPS VDD VDD P l=0.18u w=1.54u 
MM29 VDD 5 Q VDD P l=0.18u w=1.54u 
MM28 Q 5 VDD VDD P l=0.18u w=1.54u 
MM32 VDD CDN 5 VDD P l=0.184844u w=1.412u 
MM27 VDD IPS 5 VDD P l=0.184494u w=1.522u 
MM26 16 CDN VDD VDD P l=0.18u w=0.86u 
MM23 16 4 IPM VDD P l=0.18u w=0.59u 
MM25 17 2 IPM VDD P l=0.18u w=0.59u 
MM24 17 D VDD VDD P l=0.18u w=0.54u 
MM22 16 10 VDD VDD P l=0.187709u w=1.074u 
MM21 VDD 4 2 VDD P l=0.18u w=0.68u 
MM20 VDD CP 4 VDD P l=0.18u w=0.7u 
MM19 IPS 2 10 VSS N l=0.18u w=0.76u 
MM17 IPS 4 14 VSS N l=0.18u w=0.76u 
MM16 20 SDN 10 VSS N l=0.18u w=0.9u 
MM15 18 SDN 14 VSS N l=0.18u w=0.76u 
MM18 IPM 2 16 VSS N l=0.18u w=0.48u 
MM14 21 CDN 16 VSS N l=0.18u w=0.86u 
MM12 18 5 VSS VSS N l=0.18u w=0.76u 
MM11 5 IPS 19 VSS N l=0.18u w=1.07u 
MM13 VSS CDN 19 VSS N l=0.18u w=1.07u 
MM9 IPM 4 17 VSS N l=0.18u w=0.48u 
MM10 17 D VSS VSS N l=0.18u w=0.48u 
MM8 20 IPM VSS VSS N l=0.18u w=0.9u 
MM7 21 10 VSS VSS N l=0.18u w=0.86u 
MM6 VSS IPS QN VSS N l=0.18u w=1u 
MM5 VSS IPS QN VSS N l=0.18u w=1u 
MM4 VSS 5 Q VSS N l=0.18u w=1u 
MM3 VSS 5 Q VSS N l=0.18u w=1u 
MM2 VSS 4 2 VSS N l=0.18u w=0.52u 
MM1 VSS CP 4 VSS N l=0.18u w=0.52u 
.ENDS dfbrb2

.SUBCKT dfcfb1 Q QN  CDN CPN D VDD VSS
MM30 Q 2 VDD VDD P l=0.18u w=1.4u 
MM29 VDD IPS QN VDD P l=0.185306u w=1.47u 
MM26 VDD CDN 2 VDD P l=0.185652u w=1.38u 
MM24 VDD IPS 2 VDD P l=0.18u w=1.09u 
MM27 IPS 5 14 VDD P l=0.18u w=0.68u 
MM25 14 2 VDD VDD P l=0.18u w=0.68u 
MM23 IPS 7 10 VDD P l=0.18u w=0.85u 
MM28 VDD IPM 10 VDD P l=0.188008u w=1.034u 
MM22 VDD 5 7 VDD P l=0.18u w=0.68u 
MM21 VDD CPN 5 VDD P l=0.18u w=0.68u 
MM17 VDD 10 15 VDD P l=0.18u w=1.07u 
MM19 VDD CDN 15 VDD P l=0.186042u w=1.132u 
MM16 IPM 7 15 VDD P l=0.18u w=0.71u 
MM20 IPM 5 16 VDD P l=0.18u w=0.71u 
MM18 VDD D 16 VDD P l=0.18u w=0.71u 
MM13 10 5 IPS VSS N l=0.18u w=0.6u 
MM10 14 7 IPS VSS N l=0.18u w=0.59u 
MM15 10 IPM VSS VSS N l=0.18u w=0.6u 
MM14 IPM 5 15 VSS N l=0.18u w=0.48u 
MM12 15 CDN 18 VSS N l=0.18u w=0.59u 
MM9 IPM 7 16 VSS N l=0.18u w=0.48u 
MM8 14 2 VSS VSS N l=0.18u w=0.59u 
MM11 VSS CDN 17 VSS N l=0.185132u w=1.52u 
MM7 2 IPS 17 VSS N l=0.185132u w=1.52u 
MM6 VSS D 16 VSS N l=0.18u w=0.48u 
MM5 18 10 VSS VSS N l=0.18u w=0.59u 
MM4 VSS 2 Q VSS N l=0.18u w=1.06u 
MM3 QN IPS VSS VSS N l=0.186903u w=1.13u 
MM2 VSS 5 7 VSS N l=0.18u w=0.52u 
MM1 VSS CPN 5 VSS N l=0.18u w=0.52u 
.ENDS dfcfb1

.SUBCKT dfcfb2 Q QN  CDN CPN D VDD VSS
MM33 IPS 3 14 VDD P l=0.18u w=0.68u 
MM31 14 5 VDD VDD P l=0.18u w=0.68u 
MM30 Q 5 VDD VDD P l=0.185032u w=1.55u 
MM29 Q 5 VDD VDD P l=0.185623u w=1.558u 
MM32 VDD CDN 5 VDD P l=0.185652u w=1.38u 
MM27 VDD IPS 5 VDD P l=0.18u w=1.31u 
MM28 VDD IPS QN VDD P l=0.185032u w=1.55u 
MM26 QN IPS VDD VDD P l=0.18u w=1.48u 
MM25 IPS 7 9 VDD P l=0.18u w=0.85u 
MM34 VDD IPM 9 VDD P l=0.188008u w=1.034u 
MM21 VDD 9 15 VDD P l=0.18u w=1.07u 
MM23 VDD CDN 15 VDD P l=0.186042u w=1.132u 
MM20 IPM 7 15 VDD P l=0.18u w=0.71u 
MM24 IPM 3 16 VDD P l=0.18u w=0.71u 
MM22 VDD D 16 VDD P l=0.18u w=0.71u 
MM19 VDD 3 7 VDD P l=0.18u w=0.68u 
MM18 VDD CPN 3 VDD P l=0.18u w=0.68u 
MM15 9 3 IPS VSS N l=0.18u w=0.6u 
MM12 14 7 IPS VSS N l=0.18u w=0.59u 
MM17 9 IPM VSS VSS N l=0.18u w=0.6u 
MM16 IPM 3 15 VSS N l=0.18u w=0.48u 
MM14 15 CDN 18 VSS N l=0.18u w=0.59u 
MM11 IPM 7 16 VSS N l=0.18u w=0.48u 
MM10 14 5 VSS VSS N l=0.18u w=0.59u 
MM9 5 IPS 17 VSS N l=0.18u w=1.45u 
MM13 VSS CDN 17 VSS N l=0.18u w=1.45u 
MM8 VSS D 16 VSS N l=0.18u w=0.48u 
MM7 18 9 VSS VSS N l=0.18u w=0.59u 
MM6 VSS 5 Q VSS N l=0.187569u w=1.094u 
MM5 Q 5 VSS VSS N l=0.18u w=1.02u 
MM4 VSS IPS QN VSS N l=0.188235u w=1.122u 
MM3 VSS IPS QN VSS N l=0.18u w=1.04u 
MM2 VSS 3 7 VSS N l=0.18u w=0.52u 
MM1 VSS CPN 3 VSS N l=0.18u w=0.52u 
.ENDS dfcfb2

.SUBCKT dfcfq1 Q  CDN CPN D VDD VSS
MM28 VDD 2 11 VDD P l=0.18u w=1.07u 
MM26 VDD CDN 11 VDD P l=0.186042u w=1.132u 
MM24 IPM 6 11 VDD P l=0.18u w=0.71u 
MM27 IPM 3 15 VDD P l=0.18u w=0.71u 
MM25 VDD D 15 VDD P l=0.18u w=0.71u 
MM23 IPS 3 13 VDD P l=0.18u w=0.68u 
MM21 13 7 VDD VDD P l=0.18u w=0.68u 
MM22 VDD CDN 7 VDD P l=0.185652u w=1.38u 
MM19 VDD IPS 7 VDD P l=0.18u w=1.31u 
MM18 VDD 7 Q VDD P l=0.184845u w=1.61u 
MM17 IPS 6 2 VDD P l=0.18u w=0.85u 
MM20 VDD IPM 2 VDD P l=0.188008u w=1.034u 
MM16 VDD 3 6 VDD P l=0.18u w=0.68u 
MM15 VDD CPN 3 VDD P l=0.18u w=0.68u 
MM12 2 3 IPS VSS N l=0.18u w=0.6u 
MM9 13 6 IPS VSS N l=0.18u w=0.59u 
MM13 IPM 3 11 VSS N l=0.18u w=0.48u 
MM11 11 CDN 16 VSS N l=0.18u w=0.59u 
MM14 16 2 VSS VSS N l=0.18u w=0.59u 
MM8 IPM 6 15 VSS N l=0.18u w=0.48u 
MM7 13 7 VSS VSS N l=0.18u w=0.59u 
MM6 2 IPM VSS VSS N l=0.18u w=0.6u 
MM10 VSS CDN 17 VSS N l=0.185132u w=1.52u 
MM5 7 IPS 17 VSS N l=0.185132u w=1.52u 
MM4 VSS D 15 VSS N l=0.18u w=0.48u 
MM3 VSS 7 Q VSS N l=0.186903u w=1.13u 
MM2 VSS 3 6 VSS N l=0.18u w=0.52u 
MM1 VSS CPN 3 VSS N l=0.18u w=0.52u 
.ENDS dfcfq1

.SUBCKT dfcfq2 Q  CDN CPN D VDD VSS
MM26 VDD 5 11 VDD P l=0.18u w=1.07u 
MM28 VDD CDN 11 VDD P l=0.186042u w=1.132u 
MM25 IPM 6 11 VDD P l=0.18u w=0.71u 
MM29 IPM 2 15 VDD P l=0.18u w=0.71u 
MM27 VDD D 15 VDD P l=0.18u w=0.71u 
MM24 IPS 2 13 VDD P l=0.18u w=0.68u 
MM22 13 7 VDD VDD P l=0.18u w=0.68u 
MM23 VDD CDN 7 VDD P l=0.18u w=1.31u 
MM20 VDD IPS 7 VDD P l=0.185983u w=1.384u 
MM19 VDD 7 Q VDD P l=0.184845u w=1.61u 
MM18 VDD 7 Q VDD P l=0.18u w=1.54u 
MM17 IPS 6 5 VDD P l=0.18u w=0.85u 
MM21 VDD IPM 5 VDD P l=0.188008u w=1.034u 
MM16 VDD 2 6 VDD P l=0.18u w=0.68u 
MM15 VDD CPN 2 VDD P l=0.18u w=0.68u 
MM13 5 2 IPS VSS N l=0.18u w=0.6u 
MM10 13 6 IPS VSS N l=0.18u w=0.59u 
MM14 IPM 2 11 VSS N l=0.18u w=0.48u 
MM12 11 CDN 17 VSS N l=0.18u w=0.59u 
MM9 IPM 6 15 VSS N l=0.18u w=0.48u 
MM8 13 7 VSS VSS N l=0.18u w=0.59u 
MM7 5 IPM VSS VSS N l=0.18u w=0.6u 
MM11 VSS CDN 16 VSS N l=0.185132u w=1.52u 
MM6 7 IPS 16 VSS N l=0.185132u w=1.52u 
MM5 VSS D 15 VSS N l=0.18u w=0.48u 
MM4 17 5 VSS VSS N l=0.18u w=0.59u 
MM3 Q 7 VSS VSS N l=0.19717u w=1.908u 
MM2 VSS 2 6 VSS N l=0.18u w=0.52u 
MM1 VSS CPN 2 VSS N l=0.18u w=0.52u 
.ENDS dfcfq2

.SUBCKT dfcrb1 Q QN  CDN CP D VDD VSS
MM30 Q 2 VDD VDD P l=0.18u w=1.4u 
MM29 VDD IPS QN VDD P l=0.185306u w=1.47u 
MM26 VDD CDN 2 VDD P l=0.185652u w=1.38u 
MM24 VDD IPS 2 VDD P l=0.18u w=1.09u 
MM28 IPS 4 14 VDD P l=0.18u w=0.68u 
MM25 14 2 VDD VDD P l=0.18u w=0.68u 
MM23 IPS 7 10 VDD P l=0.18u w=0.85u 
MM27 VDD IPM 10 VDD P l=0.188008u w=1.034u 
MM22 VDD 7 4 VDD P l=0.18u w=0.68u 
MM21 VDD CP 7 VDD P l=0.18u w=0.68u 
MM17 VDD 10 15 VDD P l=0.18u w=1.07u 
MM20 VDD CDN 15 VDD P l=0.186042u w=1.132u 
MM18 IPM 7 15 VDD P l=0.18u w=0.71u 
MM16 IPM 4 16 VDD P l=0.18u w=0.71u 
MM19 VDD D 16 VDD P l=0.18u w=0.71u 
MM15 14 7 IPS VSS N l=0.18u w=0.59u 
MM14 10 4 IPS VSS N l=0.18u w=0.6u 
MM12 10 IPM VSS VSS N l=0.18u w=0.6u 
MM13 IPM 4 15 VSS N l=0.18u w=0.48u 
MM11 15 CDN 18 VSS N l=0.18u w=0.59u 
MM9 14 2 VSS VSS N l=0.18u w=0.59u 
MM10 VSS CDN 17 VSS N l=0.185132u w=1.52u 
MM8 2 IPS 17 VSS N l=0.185132u w=1.52u 
MM6 IPM 7 16 VSS N l=0.18u w=0.48u 
MM7 VSS D 16 VSS N l=0.18u w=0.48u 
MM5 18 10 VSS VSS N l=0.18u w=0.59u 
MM4 VSS 2 Q VSS N l=0.18u w=1.06u 
MM3 QN IPS VSS VSS N l=0.186903u w=1.13u 
MM2 VSS 7 4 VSS N l=0.18u w=0.52u 
MM1 VSS CP 7 VSS N l=0.18u w=0.52u 
.ENDS dfcrb1

.SUBCKT dfcrb2 Q QN  CDN CP D VDD VSS
MM34 IPS 2 14 VDD P l=0.18u w=0.68u 
MM31 14 5 VDD VDD P l=0.18u w=0.68u 
MM30 Q 5 VDD VDD P l=0.185032u w=1.55u 
MM29 Q 5 VDD VDD P l=0.185623u w=1.558u 
MM32 VDD CDN 5 VDD P l=0.185652u w=1.38u 
MM27 VDD IPS 5 VDD P l=0.18u w=1.31u 
MM28 VDD IPS QN VDD P l=0.185032u w=1.55u 
MM26 QN IPS VDD VDD P l=0.18u w=1.48u 
MM25 IPS 7 9 VDD P l=0.18u w=0.85u 
MM33 VDD IPM 9 VDD P l=0.188008u w=1.034u 
MM21 VDD 9 15 VDD P l=0.18u w=1.07u 
MM24 VDD CDN 15 VDD P l=0.186042u w=1.132u 
MM22 IPM 7 15 VDD P l=0.18u w=0.71u 
MM20 IPM 2 16 VDD P l=0.18u w=0.71u 
MM23 VDD D 16 VDD P l=0.18u w=0.71u 
MM19 VDD 7 2 VDD P l=0.18u w=0.68u 
MM18 VDD CP 7 VDD P l=0.18u w=0.68u 
MM17 14 7 IPS VSS N l=0.18u w=0.59u 
MM16 9 2 IPS VSS N l=0.18u w=0.6u 
MM14 9 IPM VSS VSS N l=0.18u w=0.6u 
MM15 IPM 2 15 VSS N l=0.18u w=0.48u 
MM13 15 CDN 18 VSS N l=0.18u w=0.59u 
MM11 14 5 VSS VSS N l=0.18u w=0.59u 
MM10 5 IPS 17 VSS N l=0.18u w=1.45u 
MM12 VSS CDN 17 VSS N l=0.18u w=1.45u 
MM8 IPM 7 16 VSS N l=0.18u w=0.48u 
MM9 VSS D 16 VSS N l=0.18u w=0.48u 
MM7 18 9 VSS VSS N l=0.18u w=0.59u 
MM6 VSS 5 Q VSS N l=0.187569u w=1.094u 
MM5 Q 5 VSS VSS N l=0.18u w=1.02u 
MM4 VSS IPS QN VSS N l=0.188235u w=1.122u 
MM3 VSS IPS QN VSS N l=0.18u w=1.04u 
MM2 VSS 7 2 VSS N l=0.18u w=0.52u 
MM1 VSS CP 7 VSS N l=0.18u w=0.52u 
.ENDS dfcrb2

.SUBCKT dfcrn1 QN  CDN CP D VDD VSS
MM28 VDD 2 11 VDD P l=0.18u w=1.07u 
MM27 VDD CDN 11 VDD P l=0.186042u w=1.132u 
MM25 IPM 5 11 VDD P l=0.18u w=0.71u 
MM24 IPM 6 15 VDD P l=0.18u w=0.71u 
MM26 VDD D 15 VDD P l=0.18u w=0.71u 
MM23 IPS 6 13 VDD P l=0.18u w=0.63u 
MM21 13 7 VDD VDD P l=0.18u w=0.63u 
MM20 VDD IPM 2 VDD P l=0.188008u w=1.034u 
MM17 IPS 5 2 VDD P l=0.18u w=0.8u 
MM19 VDD IPS QN VDD P l=0.184845u w=1.61u 
MM22 VDD CDN 7 VDD P l=0.185983u w=1.384u 
MM18 VDD IPS 7 VDD P l=0.18u w=1.31u 
MM16 VDD 5 6 VDD P l=0.18u w=0.68u 
MM15 VDD CP 5 VDD P l=0.18u w=0.68u 
MM14 2 6 IPS VSS N l=0.18u w=0.6u 
MM12 13 5 IPS VSS N l=0.18u w=0.59u 
MM13 IPM 6 11 VSS N l=0.18u w=0.48u 
MM10 11 CDN 16 VSS N l=0.18u w=0.59u 
MM11 16 2 VSS VSS N l=0.18u w=0.59u 
MM8 13 7 VSS VSS N l=0.18u w=0.59u 
MM7 2 IPM VSS VSS N l=0.18u w=0.6u 
MM9 VSS CDN 17 VSS N l=0.185132u w=1.52u 
MM6 7 IPS 17 VSS N l=0.185132u w=1.52u 
MM4 IPM 5 15 VSS N l=0.18u w=0.48u 
MM5 VSS D 15 VSS N l=0.18u w=0.48u 
MM3 VSS IPS QN VSS N l=0.186903u w=1.13u 
MM2 VSS 5 6 VSS N l=0.18u w=0.52u 
MM1 VSS CP 5 VSS N l=0.18u w=0.52u 
.ENDS dfcrn1

.SUBCKT dfcrn2 QN  CDN CP D VDD VSS
MM26 VDD 5 11 VDD P l=0.18u w=1.07u 
MM29 VDD CDN 11 VDD P l=0.186042u w=1.132u 
MM27 IPM 4 11 VDD P l=0.18u w=0.71u 
MM25 IPM 6 15 VDD P l=0.18u w=0.71u 
MM28 VDD D 15 VDD P l=0.18u w=0.71u 
MM24 IPS 6 13 VDD P l=0.18u w=0.63u 
MM22 13 7 VDD VDD P l=0.18u w=0.63u 
MM21 VDD IPM 5 VDD P l=0.188008u w=1.034u 
MM17 IPS 4 5 VDD P l=0.18u w=0.8u 
MM20 VDD IPS QN VDD P l=0.184845u w=1.61u 
MM19 VDD IPS QN VDD P l=0.18u w=1.54u 
MM23 VDD CDN 7 VDD P l=0.18u w=1.31u 
MM18 VDD IPS 7 VDD P l=0.185983u w=1.384u 
MM16 VDD 4 6 VDD P l=0.18u w=0.68u 
MM15 VDD CP 4 VDD P l=0.18u w=0.68u 
MM14 5 6 IPS VSS N l=0.18u w=0.6u 
MM12 13 4 IPS VSS N l=0.18u w=0.59u 
MM13 IPM 6 11 VSS N l=0.18u w=0.48u 
MM11 11 CDN 17 VSS N l=0.18u w=0.59u 
MM9 13 7 VSS VSS N l=0.18u w=0.59u 
MM8 5 IPM VSS VSS N l=0.18u w=0.6u 
MM10 VSS CDN 16 VSS N l=0.185132u w=1.52u 
MM7 7 IPS 16 VSS N l=0.185132u w=1.52u 
MM5 IPM 4 15 VSS N l=0.18u w=0.48u 
MM6 VSS D 15 VSS N l=0.18u w=0.48u 
MM4 17 5 VSS VSS N l=0.18u w=0.59u 
MM3 QN IPS VSS VSS N l=0.19717u w=1.908u 
MM2 VSS 4 6 VSS N l=0.18u w=0.52u 
MM1 VSS CP 4 VSS N l=0.18u w=0.52u 
.ENDS dfcrn2

.SUBCKT dfcrq1 Q  CDN CP D VDD VSS
MM28 VDD 2 11 VDD P l=0.18u w=1.07u 
MM27 VDD CDN 11 VDD P l=0.186042u w=1.132u 
MM25 IPM 5 11 VDD P l=0.18u w=0.71u 
MM24 IPM 6 15 VDD P l=0.18u w=0.71u 
MM26 VDD D 15 VDD P l=0.18u w=0.71u 
MM23 IPS 6 13 VDD P l=0.18u w=0.63u 
MM21 13 7 VDD VDD P l=0.18u w=0.63u 
MM20 VDD IPM 2 VDD P l=0.188008u w=1.034u 
MM17 IPS 5 2 VDD P l=0.18u w=0.8u 
MM22 VDD CDN 7 VDD P l=0.185983u w=1.384u 
MM19 VDD IPS 7 VDD P l=0.18u w=1.31u 
MM18 VDD 7 Q VDD P l=0.184845u w=1.61u 
MM16 VDD 5 6 VDD P l=0.18u w=0.68u 
MM15 VDD CP 5 VDD P l=0.18u w=0.68u 
MM14 2 6 IPS VSS N l=0.18u w=0.6u 
MM12 13 5 IPS VSS N l=0.18u w=0.59u 
MM13 IPM 6 11 VSS N l=0.18u w=0.48u 
MM10 11 CDN 16 VSS N l=0.18u w=0.59u 
MM11 16 2 VSS VSS N l=0.18u w=0.59u 
MM8 13 7 VSS VSS N l=0.18u w=0.59u 
MM7 2 IPM VSS VSS N l=0.18u w=0.6u 
MM9 VSS CDN 17 VSS N l=0.185132u w=1.52u 
MM6 7 IPS 17 VSS N l=0.185132u w=1.52u 
MM4 IPM 5 15 VSS N l=0.18u w=0.48u 
MM5 VSS D 15 VSS N l=0.18u w=0.48u 
MM3 VSS 7 Q VSS N l=0.186903u w=1.13u 
MM2 VSS 5 6 VSS N l=0.18u w=0.52u 
MM1 VSS CP 5 VSS N l=0.18u w=0.52u 
.ENDS dfcrq1

.SUBCKT dfcrq2 Q  CDN CP D VDD VSS
MM26 VDD 5 11 VDD P l=0.18u w=1.07u 
MM29 VDD CDN 11 VDD P l=0.186042u w=1.132u 
MM27 IPM 4 11 VDD P l=0.18u w=0.71u 
MM25 IPM 6 15 VDD P l=0.18u w=0.71u 
MM28 VDD D 15 VDD P l=0.18u w=0.71u 
MM24 IPS 6 13 VDD P l=0.18u w=0.63u 
MM22 13 7 VDD VDD P l=0.18u w=0.63u 
MM21 VDD IPM 5 VDD P l=0.188008u w=1.034u 
MM17 IPS 4 5 VDD P l=0.18u w=0.8u 
MM23 VDD CDN 7 VDD P l=0.18u w=1.31u 
MM20 VDD IPS 7 VDD P l=0.185983u w=1.384u 
MM19 VDD 7 Q VDD P l=0.184845u w=1.61u 
MM18 VDD 7 Q VDD P l=0.18u w=1.54u 
MM16 VDD 4 6 VDD P l=0.18u w=0.68u 
MM15 VDD CP 4 VDD P l=0.18u w=0.68u 
MM14 5 6 IPS VSS N l=0.18u w=0.6u 
MM12 13 4 IPS VSS N l=0.18u w=0.59u 
MM13 IPM 6 11 VSS N l=0.18u w=0.48u 
MM11 11 CDN 17 VSS N l=0.18u w=0.59u 
MM9 13 7 VSS VSS N l=0.18u w=0.59u 
MM8 5 IPM VSS VSS N l=0.18u w=0.6u 
MM10 VSS CDN 16 VSS N l=0.185132u w=1.52u 
MM7 7 IPS 16 VSS N l=0.185132u w=1.52u 
MM5 IPM 4 15 VSS N l=0.18u w=0.48u 
MM6 VSS D 15 VSS N l=0.18u w=0.48u 
MM4 17 5 VSS VSS N l=0.18u w=0.59u 
MM3 Q 7 VSS VSS N l=0.19717u w=1.908u 
MM2 VSS 4 6 VSS N l=0.18u w=0.52u 
MM1 VSS CP 4 VSS N l=0.18u w=0.52u 
.ENDS dfcrq2

.SUBCKT dfnfb1 Q QN  CPN D VDD VSS
MM26 8 IPM VDD VDD P l=0.18u w=1.01u 
MM25 8 3 IPS VDD P l=0.187222u w=1.08u 
MM23 IPS 4 13 VDD P l=0.18u w=0.68u 
MM24 IPM 3 14 VDD P l=0.18u w=0.6u 
MM18 VDD 8 14 VDD P l=0.18u w=0.51u 
MM21 VDD 5 13 VDD P l=0.18u w=0.44u 
MM22 IPM 4 15 VDD P l=0.18u w=0.6u 
MM19 VDD D 15 VDD P l=0.18u w=0.52u 
MM20 VDD IPS 5 VDD P l=0.18u w=0.49u 
MM17 Q 5 VDD VDD P l=0.184554u w=1.502u 
MM16 QN IPS VDD VDD P l=0.185166u w=1.51u 
MM15 VDD CPN 4 VDD P l=0.18u w=0.67u 
MM14 VDD 4 3 VDD P l=0.18u w=0.67u 
MM11 13 3 IPS VSS N l=0.18u w=0.59u 
MM8 VSS 5 13 VSS N l=0.18u w=0.43u 
MM12 IPM 3 15 VSS N l=0.18u w=0.48u 
MM10 IPM 4 14 VSS N l=0.18u w=0.48u 
MM9 IPS 4 8 VSS N l=0.18u w=0.59u 
MM13 VSS IPM 8 VSS N l=0.18u w=0.59u 
MM7 VSS IPS 5 VSS N l=0.18u w=0.46u 
MM6 VSS D 15 VSS N l=0.18u w=0.48u 
MM5 VSS 8 14 VSS N l=0.18u w=0.59u 
MM4 VSS 5 Q VSS N l=0.187091u w=1.1u 
MM3 VSS IPS QN VSS N l=0.187222u w=1.08u 
MM2 VSS CPN 4 VSS N l=0.18u w=0.52u 
MM1 VSS 4 3 VSS N l=0.18u w=0.52u 
.ENDS dfnfb1

.SUBCKT dfnfb2 Q QN  CPN D VDD VSS
MM30 7 2 IPS VDD P l=0.187222u w=1.08u 
MM28 IPS 3 13 VDD P l=0.18u w=0.68u 
MM29 IPM 2 14 VDD P l=0.18u w=0.6u 
MM23 VDD 7 14 VDD P l=0.18u w=0.51u 
MM25 VDD 5 13 VDD P l=0.18u w=0.58u 
MM27 IPM 3 15 VDD P l=0.18u w=0.6u 
MM24 VDD D 15 VDD P l=0.18u w=0.52u 
MM26 VDD IPS 5 VDD P l=0.18u w=0.59u 
MM22 7 IPM VDD VDD P l=0.18u w=1.01u 
MM21 QN IPS VDD VDD P l=0.185032u w=1.55u 
MM20 QN IPS VDD VDD P l=0.18u w=1.48u 
MM19 VDD 5 Q VDD P l=0.185032u w=1.55u 
MM18 VDD 5 Q VDD P l=0.185623u w=1.558u 
MM17 VDD CPN 3 VDD P l=0.18u w=0.67u 
MM16 VDD 3 2 VDD P l=0.18u w=0.67u 
MM14 IPS 2 13 VSS N l=0.18u w=0.59u 
MM10 VSS 5 13 VSS N l=0.18u w=0.43u 
MM15 IPM 2 15 VSS N l=0.18u w=0.48u 
MM13 IPM 3 14 VSS N l=0.18u w=0.48u 
MM12 IPS 3 7 VSS N l=0.18u w=0.59u 
MM11 VSS IPS 5 VSS N l=0.18u w=0.46u 
MM9 VSS D 15 VSS N l=0.18u w=0.48u 
MM8 VSS 7 14 VSS N l=0.18u w=0.59u 
MM7 VSS IPM 7 VSS N l=0.18u w=0.59u 
MM6 VSS IPS QN VSS N l=0.188235u w=1.122u 
MM5 VSS IPS QN VSS N l=0.18u w=1.04u 
MM4 VSS 5 Q VSS N l=0.187569u w=1.094u 
MM3 Q 5 VSS VSS N l=0.18u w=1.02u 
MM2 VSS CPN 3 VSS N l=0.18u w=0.52u 
MM1 VSS 3 2 VSS N l=0.18u w=0.52u 
.ENDS dfnfb2

.SUBCKT dfnrb1 Q QN  CP D VDD VSS
MM25 IPS 3 13 VDD P l=0.18u w=0.68u 
MM22 VDD 5 13 VDD P l=0.18u w=0.44u 
MM24 8 4 IPS VDD P l=0.187222u w=1.08u 
MM26 8 IPM VDD VDD P l=0.18u w=1.01u 
MM23 IPM 4 15 VDD P l=0.18u w=0.6u 
MM19 VDD 8 15 VDD P l=0.18u w=0.51u 
MM21 VDD IPS 5 VDD P l=0.18u w=0.49u 
MM20 VDD D 14 VDD P l=0.18u w=0.52u 
MM18 IPM 3 14 VDD P l=0.18u w=0.6u 
MM17 Q 5 VDD VDD P l=0.184554u w=1.502u 
MM16 QN IPS VDD VDD P l=0.185166u w=1.51u 
MM15 VDD 4 3 VDD P l=0.18u w=0.68u 
MM14 VDD CP 4 VDD P l=0.18u w=0.68u 
MM13 13 4 IPS VSS N l=0.18u w=0.59u 
MM8 VSS 5 13 VSS N l=0.18u w=0.43u 
MM11 IPS 3 8 VSS N l=0.18u w=0.59u 
MM12 VSS IPM 8 VSS N l=0.18u w=0.59u 
MM10 IPM 3 15 VSS N l=0.18u w=0.48u 
MM9 IPM 4 14 VSS N l=0.18u w=0.48u 
MM7 VSS IPS 5 VSS N l=0.18u w=0.46u 
MM6 VSS D 14 VSS N l=0.18u w=0.48u 
MM5 VSS 8 15 VSS N l=0.18u w=0.59u 
MM4 VSS 5 Q VSS N l=0.187222u w=1.08u 
MM3 VSS IPS QN VSS N l=0.186903u w=1.13u 
MM2 VSS 4 3 VSS N l=0.18u w=0.52u 
MM1 VSS CP 4 VSS N l=0.18u w=0.52u 
.ENDS dfnrb1

.SUBCKT dfnrb2 Q QN  CP D VDD VSS
MM30 IPS 2 13 VDD P l=0.18u w=0.68u 
MM26 VDD 5 13 VDD P l=0.18u w=0.58u 
MM29 7 3 IPS VDD P l=0.187222u w=1.08u 
MM28 IPM 3 15 VDD P l=0.18u w=0.6u 
MM24 VDD 7 15 VDD P l=0.18u w=0.51u 
MM27 VDD IPS 5 VDD P l=0.18u w=0.59u 
MM23 7 IPM VDD VDD P l=0.18u w=1.01u 
MM25 VDD D 14 VDD P l=0.18u w=0.52u 
MM22 IPM 2 14 VDD P l=0.18u w=0.6u 
MM21 QN IPS VDD VDD P l=0.185032u w=1.55u 
MM20 QN IPS VDD VDD P l=0.18u w=1.48u 
MM19 VDD 5 Q VDD P l=0.185032u w=1.55u 
MM18 VDD 5 Q VDD P l=0.185623u w=1.558u 
MM17 VDD 3 2 VDD P l=0.18u w=0.68u 
MM16 VDD CP 3 VDD P l=0.18u w=0.68u 
MM15 IPS 3 13 VSS N l=0.18u w=0.59u 
MM10 VSS 5 13 VSS N l=0.18u w=0.43u 
MM14 IPS 2 7 VSS N l=0.18u w=0.59u 
MM13 IPM 2 15 VSS N l=0.18u w=0.48u 
MM12 IPM 3 14 VSS N l=0.18u w=0.48u 
MM11 VSS IPS 5 VSS N l=0.18u w=0.46u 
MM9 VSS D 14 VSS N l=0.18u w=0.48u 
MM8 VSS 7 15 VSS N l=0.18u w=0.59u 
MM7 VSS IPM 7 VSS N l=0.18u w=0.59u 
MM6 VSS IPS QN VSS N l=0.188235u w=1.122u 
MM5 VSS IPS QN VSS N l=0.18u w=1.04u 
MM4 VSS 5 Q VSS N l=0.187569u w=1.094u 
MM3 Q 5 VSS VSS N l=0.18u w=1.02u 
MM2 VSS 3 2 VSS N l=0.18u w=0.52u 
MM1 VSS CP 3 VSS N l=0.18u w=0.52u 
.ENDS dfnrb2

.SUBCKT dfnrn1 QN  CP D VDD VSS
MM24 12 2 IPS VDD P l=0.18u w=0.68u 
MM23 7 3 IPS VDD P l=0.18u w=0.98u 
MM20 12 5 VDD VDD P l=0.18u w=0.52u 
MM22 IPM 3 14 VDD P l=0.18u w=0.6u 
MM18 VDD 7 14 VDD P l=0.18u w=0.51u 
MM21 7 IPM VDD VDD P l=0.18u w=0.98u 
MM19 VDD D 13 VDD P l=0.18u w=0.52u 
MM17 IPM 2 13 VDD P l=0.18u w=0.6u 
MM16 VDD IPS QN VDD P l=0.185166u w=1.51u 
MM15 VDD IPS 5 VDD P l=0.18u w=0.52u 
MM14 VDD 3 2 VDD P l=0.18u w=0.68u 
MM13 VDD CP 3 VDD P l=0.18u w=0.68u 
MM12 12 3 IPS VSS N l=0.18u w=0.59u 
MM7 VSS 5 12 VSS N l=0.18u w=0.43u 
MM11 IPS 2 7 VSS N l=0.18u w=0.59u 
MM10 IPM 2 14 VSS N l=0.18u w=0.48u 
MM9 IPM 3 13 VSS N l=0.18u w=0.48u 
MM8 VSS IPM 7 VSS N l=0.18u w=0.59u 
MM6 VSS D 13 VSS N l=0.18u w=0.48u 
MM5 VSS 7 14 VSS N l=0.18u w=0.59u 
MM4 5 IPS VSS VSS N l=0.18u w=0.48u 
MM3 QN IPS VSS VSS N l=0.18u w=1u 
MM2 VSS 3 2 VSS N l=0.18u w=0.52u 
MM1 VSS CP 3 VSS N l=0.18u w=0.52u 
.ENDS dfnrn1

.SUBCKT dfnrn2 QN  CP D VDD VSS
MM25 12 3 IPS VDD P l=0.18u w=0.68u 
MM24 7 4 IPS VDD P l=0.18u w=0.98u 
MM22 12 5 VDD VDD P l=0.18u w=0.52u 
MM26 7 IPM VDD VDD P l=0.18u w=0.98u 
MM23 IPM 4 14 VDD P l=0.18u w=0.6u 
MM20 VDD 7 14 VDD P l=0.18u w=0.51u 
MM21 VDD D 13 VDD P l=0.18u w=0.52u 
MM19 IPM 3 13 VDD P l=0.18u w=0.6u 
MM17 VDD IPS 5 VDD P l=0.18u w=0.52u 
MM18 VDD IPS QN VDD P l=0.185166u w=1.51u 
MM16 VDD IPS QN VDD P l=0.18u w=1.44u 
MM15 VDD 4 3 VDD P l=0.18u w=0.68u 
MM14 VDD CP 4 VDD P l=0.18u w=0.68u 
MM13 12 4 IPS VSS N l=0.18u w=0.59u 
MM8 VSS 5 12 VSS N l=0.18u w=0.43u 
MM11 IPS 3 7 VSS N l=0.18u w=0.59u 
MM12 VSS IPM 7 VSS N l=0.18u w=0.59u 
MM10 IPM 3 14 VSS N l=0.18u w=0.48u 
MM9 IPM 4 13 VSS N l=0.18u w=0.48u 
MM7 VSS D 13 VSS N l=0.18u w=0.48u 
MM6 VSS 7 14 VSS N l=0.18u w=0.59u 
MM4 VSS IPS 5 VSS N l=0.18u w=0.48u 
MM5 QN IPS VSS VSS N l=0.188385u w=1.102u 
MM3 QN IPS VSS VSS N l=0.18u w=1.02u 
MM2 VSS 4 3 VSS N l=0.18u w=0.52u 
MM1 VSS CP 4 VSS N l=0.18u w=0.52u 
.ENDS dfnrn2

.SUBCKT dfnrq1 Q  CP D VDD VSS
MM24 12 2 IPS VDD P l=0.18u w=0.68u 
MM23 7 3 IPS VDD P l=0.18u w=0.98u 
MM20 12 5 VDD VDD P l=0.18u w=0.52u 
MM22 IPM 3 14 VDD P l=0.18u w=0.6u 
MM18 VDD 7 14 VDD P l=0.18u w=0.51u 
MM21 7 IPM VDD VDD P l=0.18u w=0.98u 
MM19 VDD D 13 VDD P l=0.18u w=0.52u 
MM17 IPM 2 13 VDD P l=0.18u w=0.6u 
MM16 VDD IPS 5 VDD P l=0.18u w=0.52u 
MM15 VDD 5 Q VDD P l=0.185166u w=1.51u 
MM14 VDD 3 2 VDD P l=0.18u w=0.68u 
MM13 VDD CP 3 VDD P l=0.18u w=0.68u 
MM12 12 3 IPS VSS N l=0.18u w=0.59u 
MM7 VSS 5 12 VSS N l=0.18u w=0.43u 
MM11 IPS 2 7 VSS N l=0.18u w=0.59u 
MM10 IPM 2 14 VSS N l=0.18u w=0.48u 
MM9 IPM 3 13 VSS N l=0.18u w=0.48u 
MM8 VSS IPM 7 VSS N l=0.18u w=0.59u 
MM6 VSS D 13 VSS N l=0.18u w=0.48u 
MM5 VSS 7 14 VSS N l=0.18u w=0.59u 
MM4 VSS IPS 5 VSS N l=0.18u w=0.48u 
MM3 Q 5 VSS VSS N l=0.18u w=1u 
MM2 VSS 3 2 VSS N l=0.18u w=0.52u 
MM1 VSS CP 3 VSS N l=0.18u w=0.52u 
.ENDS dfnrq1

.SUBCKT dfnrq2 Q  CP D VDD VSS
MM25 12 3 IPS VDD P l=0.18u w=0.68u 
MM24 7 4 IPS VDD P l=0.18u w=0.98u 
MM22 12 5 VDD VDD P l=0.18u w=0.52u 
MM26 7 IPM VDD VDD P l=0.18u w=0.98u 
MM23 IPM 4 14 VDD P l=0.18u w=0.6u 
MM20 VDD 7 14 VDD P l=0.18u w=0.51u 
MM21 VDD D 13 VDD P l=0.18u w=0.52u 
MM19 IPM 3 13 VDD P l=0.18u w=0.6u 
MM18 VDD IPS 5 VDD P l=0.18u w=0.51u 
MM17 VDD 5 Q VDD P l=0.1852u w=1.5u 
MM16 VDD 5 Q VDD P l=0.18u w=1.43u 
MM15 VDD 4 3 VDD P l=0.18u w=0.68u 
MM14 VDD CP 4 VDD P l=0.18u w=0.68u 
MM13 12 4 IPS VSS N l=0.18u w=0.59u 
MM8 VSS 5 12 VSS N l=0.18u w=0.43u 
MM11 IPS 3 7 VSS N l=0.18u w=0.59u 
MM12 VSS IPM 7 VSS N l=0.18u w=0.59u 
MM10 IPM 3 14 VSS N l=0.18u w=0.48u 
MM9 IPM 4 13 VSS N l=0.18u w=0.48u 
MM7 VSS D 13 VSS N l=0.18u w=0.48u 
MM6 VSS 7 14 VSS N l=0.18u w=0.59u 
MM5 VSS IPS 5 VSS N l=0.18u w=0.48u 
MM4 Q 5 VSS VSS N l=0.187569u w=1.094u 
MM3 Q 5 VSS VSS N l=0.18u w=1.02u 
MM2 VSS 4 3 VSS N l=0.18u w=0.52u 
MM1 VSS CP 4 VSS N l=0.18u w=0.52u 
.ENDS dfnrq2

.SUBCKT dfpfb1 Q QN  CPN D SDN VDD VSS
MM30 14 SDN VDD VDD P l=0.186207u w=1.102u 
MM28 14 3 IPS VDD P l=0.18u w=0.81u 
MM29 VDD SDN 9 VDD P l=0.18u w=0.78u 
MM25 9 6 IPS VDD P l=0.18u w=0.63u 
MM27 14 4 VDD VDD P l=0.18u w=1.11u 
MM26 9 IPM VDD VDD P l=0.187884u w=1.271u 
MM24 4 IPS VDD VDD P l=0.18u w=1.25u 
MM23 15 3 IPM VDD P l=0.18u w=0.59u 
MM22 VDD D 15 VDD P l=0.18u w=0.59u 
MM21 VDD 9 16 VDD P l=0.18u w=0.51u 
MM20 IPM 6 16 VDD P l=0.18u w=0.59u 
MM19 Q 4 VDD VDD P l=0.18u w=1.4u 
MM18 QN IPS VDD VDD P l=0.185306u w=1.47u 
MM17 VDD 3 6 VDD P l=0.18u w=0.65u 
MM16 VDD CPN 3 VDD P l=0.18u w=0.7u 
MM15 18 SDN 9 VSS N l=0.18u w=0.99u 
MM12 IPS 3 9 VSS N l=0.18u w=0.71u 
MM11 IPM 6 15 VSS N l=0.18u w=1.12u 
MM7 15 D VSS VSS N l=0.18u w=0.48u 
MM13 IPM 3 16 VSS N l=0.188274u w=1.211u 
MM14 14 SDN 17 VSS N l=0.18u w=0.71u 
MM10 IPS 6 14 VSS N l=0.18u w=0.71u 
MM9 17 4 VSS VSS N l=0.18u w=0.71u 
MM8 4 IPS VSS VSS N l=0.18u w=0.68u 
MM6 16 9 VSS VSS N l=0.18u w=0.54u 
MM5 18 IPM VSS VSS N l=0.18u w=0.99u 
MM4 VSS 4 Q VSS N l=0.18u w=1.06u 
MM3 VSS IPS QN VSS N l=0.186903u w=1.13u 
MM2 VSS 3 6 VSS N l=0.18u w=0.52u 
MM1 VSS CPN 3 VSS N l=0.18u w=0.52u 
.ENDS dfpfb1

.SUBCKT dfpfb2 Q QN  CPN D SDN VDD VSS
MM34 14 SDN VDD VDD P l=0.186207u w=1.102u 
MM32 14 3 IPS VDD P l=0.18u w=0.81u 
MM33 VDD SDN 9 VDD P l=0.18u w=0.78u 
MM31 9 4 IPS VDD P l=0.18u w=0.63u 
MM30 14 5 VDD VDD P l=0.18u w=1.11u 
MM29 9 IPM VDD VDD P l=0.187884u w=1.271u 
MM28 VDD 5 Q VDD P l=0.185032u w=1.55u 
MM27 VDD 5 Q VDD P l=0.185623u w=1.558u 
MM25 5 IPS VDD VDD P l=0.18u w=1.25u 
MM26 QN IPS VDD VDD P l=0.185032u w=1.55u 
MM24 VDD IPS QN VDD P l=0.18u w=1.48u 
MM23 15 3 IPM VDD P l=0.18u w=0.59u 
MM22 VDD D 15 VDD P l=0.18u w=0.59u 
MM21 VDD 9 16 VDD P l=0.18u w=0.51u 
MM20 IPM 4 16 VDD P l=0.18u w=0.59u 
MM19 VDD 3 4 VDD P l=0.18u w=0.65u 
MM18 VDD CPN 3 VDD P l=0.18u w=0.7u 
MM17 18 SDN 9 VSS N l=0.18u w=0.99u 
MM14 IPS 3 9 VSS N l=0.18u w=0.71u 
MM13 IPM 4 15 VSS N l=0.18u w=1.12u 
MM9 15 D VSS VSS N l=0.18u w=0.48u 
MM15 IPM 3 16 VSS N l=0.188274u w=1.211u 
MM16 14 SDN 17 VSS N l=0.18u w=0.71u 
MM12 IPS 4 14 VSS N l=0.18u w=0.71u 
MM11 17 5 VSS VSS N l=0.18u w=0.71u 
MM10 5 IPS VSS VSS N l=0.18u w=0.68u 
MM8 16 9 VSS VSS N l=0.18u w=0.54u 
MM7 18 IPM VSS VSS N l=0.18u w=0.99u 
MM6 Q 5 VSS VSS N l=0.187569u w=1.094u 
MM5 Q 5 VSS VSS N l=0.18u w=1.02u 
MM4 QN IPS VSS VSS N l=0.188235u w=1.122u 
MM3 QN IPS VSS VSS N l=0.18u w=1.04u 
MM2 VSS 3 4 VSS N l=0.18u w=0.52u 
MM1 VSS CPN 3 VSS N l=0.18u w=0.52u 
.ENDS dfpfb2

.SUBCKT dfprb1 Q QN  CP D SDN VDD VSS
MM30 14 2 IPS VDD P l=0.18u w=0.81u 
MM25 8 6 IPS VDD P l=0.18u w=0.63u 
MM29 14 SDN VDD VDD P l=0.186207u w=1.102u 
MM28 VDD SDN 8 VDD P l=0.18u w=0.78u 
MM27 14 4 VDD VDD P l=0.18u w=1.11u 
MM26 8 IPM VDD VDD P l=0.187884u w=1.271u 
MM24 4 IPS VDD VDD P l=0.18u w=1.25u 
MM22 VDD 8 16 VDD P l=0.18u w=0.51u 
MM20 16 6 IPM VDD P l=0.18u w=0.59u 
MM23 15 2 IPM VDD P l=0.18u w=0.59u 
MM21 VDD D 15 VDD P l=0.18u w=0.59u 
MM19 Q 4 VDD VDD P l=0.18u w=1.4u 
MM18 QN IPS VDD VDD P l=0.185306u w=1.47u 
MM17 VDD CP 6 VDD P l=0.18u w=0.7u 
MM16 VDD 6 2 VDD P l=0.18u w=0.65u 
MM14 IPS 2 8 VSS N l=0.18u w=0.71u 
MM13 18 SDN 8 VSS N l=0.18u w=0.99u 
MM11 IPM 6 15 VSS N l=0.18u w=1.12u 
MM6 15 D VSS VSS N l=0.18u w=0.48u 
MM15 IPM 2 16 VSS N l=0.188274u w=1.211u 
MM12 14 SDN 17 VSS N l=0.18u w=0.71u 
MM10 IPS 6 14 VSS N l=0.18u w=0.71u 
MM9 17 4 VSS VSS N l=0.18u w=0.71u 
MM8 4 IPS VSS VSS N l=0.18u w=0.68u 
MM7 16 8 VSS VSS N l=0.18u w=0.54u 
MM5 18 IPM VSS VSS N l=0.18u w=0.99u 
MM4 VSS 4 Q VSS N l=0.18u w=1.06u 
MM3 VSS IPS QN VSS N l=0.186903u w=1.13u 
MM2 VSS CP 6 VSS N l=0.18u w=0.52u 
MM1 VSS 6 2 VSS N l=0.18u w=0.52u 
.ENDS dfprb1

.SUBCKT dfprb2 Q QN  CP D SDN VDD VSS
MM34 14 2 IPS VDD P l=0.18u w=0.81u 
MM31 8 4 IPS VDD P l=0.18u w=0.63u 
MM33 14 SDN VDD VDD P l=0.186207u w=1.102u 
MM32 VDD SDN 8 VDD P l=0.18u w=0.78u 
MM30 14 5 VDD VDD P l=0.18u w=1.11u 
MM29 8 IPM VDD VDD P l=0.187884u w=1.271u 
MM28 VDD 5 Q VDD P l=0.185032u w=1.55u 
MM27 VDD 5 Q VDD P l=0.185623u w=1.558u 
MM25 5 IPS VDD VDD P l=0.18u w=1.25u 
MM26 QN IPS VDD VDD P l=0.185032u w=1.55u 
MM24 VDD IPS QN VDD P l=0.18u w=1.48u 
MM22 VDD 8 16 VDD P l=0.18u w=0.51u 
MM20 16 4 IPM VDD P l=0.18u w=0.59u 
MM23 15 2 IPM VDD P l=0.18u w=0.59u 
MM21 VDD D 15 VDD P l=0.18u w=0.59u 
MM19 VDD CP 4 VDD P l=0.18u w=0.7u 
MM18 VDD 4 2 VDD P l=0.18u w=0.65u 
MM16 IPS 2 8 VSS N l=0.18u w=0.71u 
MM15 18 SDN 8 VSS N l=0.18u w=0.99u 
MM13 IPM 4 15 VSS N l=0.18u w=1.12u 
MM8 15 D VSS VSS N l=0.18u w=0.48u 
MM17 IPM 2 16 VSS N l=0.188274u w=1.211u 
MM14 14 SDN 17 VSS N l=0.18u w=0.71u 
MM12 IPS 4 14 VSS N l=0.18u w=0.71u 
MM11 17 5 VSS VSS N l=0.18u w=0.71u 
MM10 5 IPS VSS VSS N l=0.18u w=0.68u 
MM9 16 8 VSS VSS N l=0.18u w=0.54u 
MM7 18 IPM VSS VSS N l=0.18u w=0.99u 
MM6 Q 5 VSS VSS N l=0.187569u w=1.094u 
MM5 Q 5 VSS VSS N l=0.18u w=1.02u 
MM4 QN IPS VSS VSS N l=0.188235u w=1.122u 
MM3 QN IPS VSS VSS N l=0.18u w=1.04u 
MM2 VSS CP 4 VSS N l=0.18u w=0.52u 
MM1 VSS 4 2 VSS N l=0.18u w=0.52u 
.ENDS dfprb2

.SUBCKT dl01d1 Z  I VDD VSS
MM8 VDD 2 4 VDD P l=0.38u w=0.42u 
MM7 VDD I 2 VDD P l=0.184875u w=1.6u 
MM6 VDD 4 5 VDD P l=0.4u w=0.42u 
MM5 VDD 5 Z VDD P l=0.18u w=1.48u 
MM4 5 4 VSS VSS N l=0.7u w=0.45u 
MM3 Z 5 VSS VSS N l=0.18u w=0.46u 
MM2 VSS 2 4 VSS N l=0.4u w=0.47u 
MM1 2 I VSS VSS N l=0.18u w=0.42u 
.ENDS dl01d1

.SUBCKT dl02d1 Z  I VDD VSS
MM8 VDD 2 4 VDD P l=0.8u w=0.42u 
MM7 VDD I 2 VDD P l=0.184875u w=1.6u 
MM6 VDD 4 5 VDD P l=0.89u w=0.42u 
MM5 VDD 5 Z VDD P l=0.18u w=1.48u 
MM4 VSS 4 5 VSS N l=0.85u w=0.45u 
MM3 VSS 5 Z VSS N l=0.18u w=0.46u 
MM2 VSS 2 4 VSS N l=1.1u w=0.47u 
MM1 2 I VSS VSS N l=0.18u w=0.42u 
.ENDS dl02d1

.SUBCKT dl03d1 Z  I VDD VSS
MM8 VDD 2 5 VDD P l=1.32u w=0.48u 
MM7 VDD I 2 VDD P l=0.184875u w=1.6u 
MM6 Z 4 VDD VDD P l=0.184756u w=1.64u 
MM5 VDD 5 4 VDD P l=1.9u w=0.42u 
MM4 Z 4 VSS VSS N l=0.18u w=0.42u 
MM3 4 5 VSS VSS N l=1.5u w=0.45u 
MM2 VSS 2 5 VSS N l=1.25u w=0.47u 
MM1 2 I VSS VSS N l=0.18u w=0.42u 
.ENDS dl03d1

.SUBCKT dl04d1 Z  I VDD VSS
MM8 VDD 2 5 VDD P l=2.1u w=0.48u 
MM7 VDD I 2 VDD P l=0.184875u w=1.6u 
MM6 Z 4 VDD VDD P l=0.184756u w=1.64u 
MM5 VDD 5 4 VDD P l=3.65u w=0.42u 
MM4 VSS 4 Z VSS N l=0.18u w=0.42u 
MM3 VSS 5 4 VSS N l=1.71u w=0.45u 
MM2 5 2 VSS VSS N l=2.54u w=0.42u 
MM1 2 I VSS VSS N l=0.18u w=0.42u 
.ENDS dl04d1

.SUBCKT feedth  VDD VSS

.ENDS feedth

.SUBCKT feedth3  VDD VSS

.ENDS feedth3

.SUBCKT feedth9  VDD VSS

.ENDS feedth9

.SUBCKT inv0d0 ZN  I VDD VSS
MM2 VDD I ZN VDD P l=0.18u w=0.36u 
MM1 ZN I VSS VSS N l=0.18u w=0.24u 
.ENDS inv0d0

.SUBCKT inv0d1 ZN  I VDD VSS
MM2 ZN I VDD VDD P l=0.18u w=1.48u 
MM1 VSS I ZN VSS N l=0.18u w=1.01u 
.ENDS inv0d1

.SUBCKT inv0d2 ZN  I VDD VSS
MM4 ZN I VDD VDD P l=0.184436u w=1.542u 
MM3 ZN I VDD VDD P l=0.18u w=1.48u 
MM2 VSS I ZN VSS N l=0.185937u w=1.152u 
MM1 VSS I ZN VSS N l=0.18u w=1.09u 
.ENDS inv0d2

.SUBCKT inv0d4 ZN  I VDD VSS
MM8 ZN I VDD VDD P l=0.184436u w=1.542u 
MM7 ZN I VDD VDD P l=0.18u w=1.48u 
MM6 ZN I VDD VDD P l=0.18u w=1.48u 
MM5 VDD I ZN VDD P l=0.184436u w=1.542u 
MM4 VSS I ZN VSS N l=0.185937u w=1.152u 
MM2 VSS I ZN VSS N l=0.18u w=1.09u 
MM3 ZN I VSS VSS N l=0.185937u w=1.152u 
MM1 ZN I VSS VSS N l=0.18u w=1.09u 
.ENDS inv0d4

.SUBCKT inv0d7 ZN  I VDD VSS
MM9 VDD I ZN VDD P l=0.183786u w=2.06u 
MM8 VDD I ZN VDD P l=0.18u w=1.99u 
MM7 ZN I VDD VDD P l=0.183786u w=2.06u 
MM6 ZN I VDD VDD P l=0.18u w=1.99u 
MM5 VDD I ZN VDD P l=0.183786u w=2.06u 
MM3 VSS I ZN VSS N l=0.184091u w=1.672u 
MM2 VSS I ZN VSS N l=0.18u w=1.61u 
MM4 VSS I ZN VSS N l=0.185461u w=1.692u 
MM1 VSS I ZN VSS N l=0.18u w=1.61u 
.ENDS inv0d7

.SUBCKT inv0da ZN  I VDD VSS
MM13 ZN I VDD VDD P l=0.183786u w=2.06u 
MM12 VDD I ZN VDD P l=0.185065u w=1.54u 
MM11 ZN I VDD VDD P l=0.183786u w=2.06u 
MM10 ZN I VDD VDD P l=0.183786u w=2.06u 
MM9 VDD I ZN VDD P l=0.183786u w=2.06u 
MM8 VDD I ZN VDD P l=0.183786u w=2.06u 
MM7 ZN I VDD VDD P l=0.183786u w=2.06u 
MM6 VSS I ZN VSS N l=0.184091u w=1.672u 
MM3 VSS I ZN VSS N l=0.18u w=1.61u 
MM5 VSS I ZN VSS N l=0.184091u w=1.672u 
MM2 ZN I VSS VSS N l=0.18u w=1.61u 
MM4 VSS I ZN VSS N l=0.184091u w=1.672u 
MM1 VSS I ZN VSS N l=0.18u w=1.61u 
.ENDS inv0da

.SUBCKT invbd2 ZN  I VDD VSS
MM5 VDD I ZN VDD P l=0.189901u w=1.624u 
MM4 ZN I VDD VDD P l=0.185032u w=1.55u 
MM3 ZN I VDD VDD P l=0.185032u w=1.55u 
MM2 ZN I VSS VSS N l=0.18u w=0.8u 
MM1 ZN I VSS VSS N l=0.18u w=0.8u 
.ENDS invbd2

.SUBCKT invbd4 ZN  I VDD VSS
MM7 VDD I ZN VDD P l=0.184021u w=1.94u 
MM6 VDD I ZN VDD P l=0.184259u w=1.944u 
MM5 VDD I ZN VDD P l=0.18u w=1.87u 
MM4 VDD I ZN VDD P l=0.184259u w=1.944u 
MM3 ZN I VDD VDD P l=0.187116u w=1.366u 
MM2 VSS I ZN VSS N l=0.193262u w=1.692u 
MM1 VSS I ZN VSS N l=0.193341u w=1.682u 
.ENDS invbd4

.SUBCKT invtd1 ZN  EN I VDD VSS
MM5 4 EN VDD VDD P l=0.18u w=0.95u 
MM6 8 EN VDD VDD P l=0.184497u w=1.948u 
MM4 8 I ZN VDD P l=0.18u w=1.87u 
MM3 4 EN VSS VSS N l=0.18u w=0.63u 
MM2 VSS 4 7 VSS N l=0.184914u w=1.392u 
MM1 7 I ZN VSS N l=0.18u w=1.33u 
.ENDS invtd1

.SUBCKT invtd2 ZN  EN I VDD VSS
MM8 4 EN VDD VDD P l=0.18u w=0.95u 
MM10 ZN EN 9 VDD P l=0.187856u w=1.581u 
MM7 VDD I 9 VDD P l=0.187856u w=1.581u 
MM9 10 EN VDD VDD P l=0.185659u w=1.548u 
MM6 ZN I 10 VDD P l=0.18u w=1.47u 
MM5 4 EN VSS VSS N l=0.18u w=0.63u 
MM3 7 4 VSS VSS N l=0.188802u w=1.411u 
MM2 7 I ZN VSS N l=0.188802u w=1.411u 
MM1 8 I ZN VSS N l=0.18u w=1.26u 
MM4 VSS 4 8 VSS N l=0.185174u w=1.322u 
.ENDS invtd2

.SUBCKT invtd4 ZN  EN I VDD VSS
MM16 VDD 2 4 VDD P l=0.18u w=1.48u 
MM15 VDD I 2 VDD P l=0.18u w=0.6u 
MM13 ZN 4 VDD VDD P l=0.189036u w=1.514u 
MM14 VDD 4 ZN VDD P l=0.185656u w=1.464u 
MM12 VDD 4 ZN VDD P l=0.18u w=1.39u 
MM11 VDD 5 4 VDD P l=0.18u w=1.06u 
MM10 7 EN 4 VDD P l=0.18u w=1.12u 
MM9 5 EN VDD VDD P l=0.18u w=0.6u 
MM8 VSS 2 7 VSS N l=0.18u w=1.04u 
MM6 ZN 7 VSS VSS N l=0.18607u w=1.364u 
MM7 ZN 7 VSS VSS N l=0.18607u w=1.364u 
MM5 ZN 7 VSS VSS N l=0.18u w=1.29u 
MM4 VSS I 2 VSS N l=0.18u w=0.44u 
MM3 4 5 7 VSS N l=0.186656u w=1.244u 
MM2 VSS EN 7 VSS N l=0.185552u w=1.232u 
MM1 VSS EN 5 VSS N l=0.18u w=0.54u 
.ENDS invtd4

.SUBCKT invtd7 ZN  EN I VDD VSS
MM22 3 2 VDD VDD P l=0.18u w=1.48u 
MM21 ZN 3 VDD VDD P l=0.185656u w=1.464u 
MM20 ZN 3 VDD VDD P l=0.18u w=1.39u 
MM19 VDD 3 ZN VDD P l=0.18u w=1.39u 
MM18 VDD 3 ZN VDD P l=0.185656u w=1.464u 
MM17 VDD 3 ZN VDD P l=0.18u w=1.39u 
MM16 VDD 3 ZN VDD P l=0.185656u w=1.464u 
MM15 2 I VDD VDD P l=0.18u w=0.6u 
MM14 VDD 5 3 VDD P l=0.18u w=1.06u 
MM13 7 EN 3 VDD P l=0.18u w=1.12u 
MM12 5 EN VDD VDD P l=0.18u w=0.6u 
MM11 VSS 2 7 VSS N l=0.18u w=1.04u 
MM9 ZN 7 VSS VSS N l=0.186115u w=1.354u 
MM7 VSS 7 ZN VSS N l=0.18u w=1.28u 
MM8 ZN 7 VSS VSS N l=0.186115u w=1.354u 
MM6 ZN 7 VSS VSS N l=0.18u w=1.28u 
MM10 VSS 7 ZN VSS N l=0.186115u w=1.354u 
MM5 VSS 7 ZN VSS N l=0.18u w=1.28u 
MM4 VSS I 2 VSS N l=0.18u w=0.44u 
MM3 3 5 7 VSS N l=0.186656u w=1.244u 
MM2 VSS EN 7 VSS N l=0.185552u w=1.232u 
MM1 VSS EN 5 VSS N l=0.18u w=0.54u 
.ENDS invtd7

.SUBCKT invtda ZN  EN I VDD VSS
MM26 VDD 2 3 VDD P l=0.18u w=1.34u 
MM25 ZN 3 VDD VDD P l=0.185656u w=1.464u 
MM24 VDD 3 ZN VDD P l=0.18u w=1.39u 
MM23 ZN 3 VDD VDD P l=0.18u w=1.39u 
MM22 ZN 3 VDD VDD P l=0.185656u w=1.464u 
MM21 ZN 3 VDD VDD P l=0.18u w=1.39u 
MM20 VDD 3 ZN VDD P l=0.185656u w=1.464u 
MM19 ZN 3 VDD VDD P l=0.18u w=1.39u 
MM18 ZN 3 VDD VDD P l=0.185656u w=1.464u 
MM17 2 I VDD VDD P l=0.18u w=0.6u 
MM15 7 EN 3 VDD P l=0.18u w=1.05u 
MM16 VDD 5 3 VDD P l=0.18u w=1.05u 
MM14 5 EN VDD VDD P l=0.18u w=0.6u 
MM13 VSS 2 7 VSS N l=0.187113u w=1.164u 
MM11 ZN 7 VSS VSS N l=0.186115u w=1.354u 
MM8 VSS 7 ZN VSS N l=0.18u w=1.28u 
MM10 VSS 7 ZN VSS N l=0.186115u w=1.354u 
MM7 ZN 7 VSS VSS N l=0.18u w=1.28u 
MM9 VSS 7 ZN VSS N l=0.186115u w=1.354u 
MM6 VSS 7 ZN VSS N l=0.18u w=1.28u 
MM12 ZN 7 VSS VSS N l=0.186115u w=1.354u 
MM5 ZN 7 VSS VSS N l=0.18u w=1.28u 
MM4 VSS I 2 VSS N l=0.18u w=0.44u 
MM3 3 5 7 VSS N l=0.186656u w=1.244u 
MM2 VSS EN 7 VSS N l=0.185552u w=1.232u 
MM1 VSS EN 5 VSS N l=0.18u w=0.54u 
.ENDS invtda

.SUBCKT jkbrb1 Q QN  CDN CP J KZ SDN VDD VSS
MM42 VDD CP 3 VDD P l=0.18u w=0.64u 
MM41 VDD 3 8 VDD P l=0.18u w=0.65u 
MM40 VDD SDN 11 VDD P l=0.18u w=0.54u 
MM38 VDD 6 11 VDD P l=0.18u w=0.69u 
MM39 6 CDN VDD VDD P l=0.18607u w=1.364u 
MM37 6 IPS VDD VDD P l=0.18u w=1.29u 
MM36 20 3 IPM VDD P l=0.18u w=0.6u 
MM35 IPM 8 19 VDD P l=0.18u w=0.6u 
MM34 26 KZ 19 VDD P l=0.18u w=0.92u 
MM33 25 J 19 VDD P l=0.18u w=0.92u 
MM32 25 11 VDD VDD P l=0.18u w=0.92u 
MM31 26 12 VDD VDD P l=0.18u w=0.92u 
MM30 Q 6 VDD VDD P l=0.18u w=1.43u 
MM29 QN IPS VDD VDD P l=0.18u w=1.43u 
MM28 IPS 3 13 VDD P l=0.18u w=0.94u 
MM27 IPS 8 11 VDD P l=0.18u w=0.59u 
MM25 VDD CDN 20 VDD P l=0.18u w=0.72u 
MM24 VDD 13 20 VDD P l=0.18u w=0.72u 
MM26 13 SDN VDD VDD P l=0.18u w=0.86u 
MM23 VDD IPM 13 VDD P l=0.18u w=0.86u 
MM22 12 11 VDD VDD P l=0.18u w=0.5u 
MM21 IPS 3 11 VSS N l=0.18u w=0.66u 
MM20 13 8 IPS VSS N l=0.18u w=0.66u 
MM19 21 SDN 11 VSS N l=0.18u w=0.66u 
MM17 21 6 VSS VSS N l=0.18u w=0.66u 
MM16 6 IPS 22 VSS N l=0.18u w=1.05u 
MM18 22 CDN VSS VSS N l=0.18u w=1.05u 
MM10 19 12 18 VSS N l=0.18u w=0.72u 
MM14 20 8 IPM VSS N l=0.18u w=0.88u 
MM15 19 3 IPM VSS N l=0.18u w=0.88u 
MM13 19 KZ 18 VSS N l=0.18u w=0.88u 
MM11 18 11 VSS VSS N l=0.18u w=0.88u 
MM12 18 J VSS VSS N l=0.18u w=0.72u 
MM9 VSS 6 Q VSS N l=0.18u w=0.95u 
MM8 VSS IPS QN VSS N l=0.18u w=0.95u 
MM7 3 CP VSS VSS N l=0.18u w=0.54u 
MM6 8 3 VSS VSS N l=0.18u w=0.54u 
MM5 24 SDN 13 VSS N l=0.18u w=0.99u 
MM4 VSS CDN 23 VSS N l=0.18u w=0.68u 
MM3 23 13 20 VSS N l=0.18u w=0.68u 
MM2 VSS IPM 24 VSS N l=0.18u w=0.99u 
MM1 VSS 11 12 VSS N l=0.18u w=0.48u 
.ENDS jkbrb1

.SUBCKT jkbrb2 Q QN  CDN CP J KZ SDN VDD VSS
MM46 VDD CP 3 VDD P l=0.18u w=0.64u 
MM45 VDD 3 8 VDD P l=0.18u w=0.65u 
MM44 11 SDN VDD VDD P l=0.18u w=0.54u 
MM39 11 7 VDD VDD P l=0.18u w=0.69u 
MM43 7 CDN VDD VDD P l=0.18u w=1.47u 
MM42 7 IPS VDD VDD P l=0.185363u w=1.544u 
MM41 QN IPS VDD VDD P l=0.185505u w=1.504u 
MM40 QN IPS VDD VDD P l=0.18u w=1.43u 
MM38 Q 7 VDD VDD P l=0.185505u w=1.504u 
MM37 Q 7 VDD VDD P l=0.18u w=1.43u 
MM36 20 3 IPM VDD P l=0.18u w=0.6u 
MM35 IPM 8 19 VDD P l=0.18u w=0.6u 
MM34 26 KZ 19 VDD P l=0.18u w=0.92u 
MM33 25 J 19 VDD P l=0.18u w=0.92u 
MM32 25 11 VDD VDD P l=0.18u w=0.92u 
MM31 26 12 VDD VDD P l=0.18u w=0.92u 
MM30 IPS 3 13 VDD P l=0.18u w=0.94u 
MM29 IPS 8 11 VDD P l=0.18u w=0.59u 
MM27 VDD CDN 20 VDD P l=0.18u w=0.72u 
MM26 VDD 13 20 VDD P l=0.18u w=0.72u 
MM28 13 SDN VDD VDD P l=0.18u w=0.86u 
MM25 VDD IPM 13 VDD P l=0.18u w=0.86u 
MM24 12 11 VDD VDD P l=0.18u w=0.5u 
MM23 3 CP VSS VSS N l=0.18u w=0.54u 
MM22 8 3 VSS VSS N l=0.18u w=0.54u 
MM21 11 3 IPS VSS N l=0.18u w=0.66u 
MM20 IPS 8 13 VSS N l=0.18u w=0.66u 
MM19 11 SDN 22 VSS N l=0.18u w=0.66u 
MM17 7 IPS 21 VSS N l=0.18u w=1.08u 
MM18 21 CDN VSS VSS N l=0.18u w=1.08u 
MM16 VSS 7 22 VSS N l=0.18u w=0.66u 
MM10 19 12 18 VSS N l=0.18u w=0.72u 
MM14 20 8 IPM VSS N l=0.18u w=0.88u 
MM15 19 3 IPM VSS N l=0.18u w=0.88u 
MM13 19 KZ 18 VSS N l=0.18u w=0.88u 
MM11 18 11 VSS VSS N l=0.18u w=0.88u 
MM12 18 J VSS VSS N l=0.18u w=0.72u 
MM9 VSS IPS QN VSS N l=0.186603u w=1.254u 
MM8 VSS IPS QN VSS N l=0.18u w=1.18u 
MM7 VSS 7 Q VSS N l=0.186603u w=1.254u 
MM6 Q 7 VSS VSS N l=0.18u w=1.18u 
MM5 24 SDN 13 VSS N l=0.18u w=0.99u 
MM4 VSS CDN 23 VSS N l=0.18u w=0.68u 
MM3 23 13 20 VSS N l=0.18u w=0.68u 
MM2 VSS IPM 24 VSS N l=0.18u w=0.99u 
MM1 VSS 11 12 VSS N l=0.18u w=0.48u 
.ENDS jkbrb2

.SUBCKT labhb1 Q QN  CDN D E SDN VDD VSS
MM28 VDD 2 6 VDD P l=0.18u w=0.57u 
MM27 VDD 2 8 VDD P l=0.18u w=0.77u 
MM26 8 3 IPM VDD P l=0.18u w=0.67u 
MM25 16 4 IPM VDD P l=0.18u w=0.72u 
MM24 VDD CDN 8 VDD P l=0.186628u w=1.032u 
MM23 VDD 6 Q VDD P l=0.186497u w=1.496u 
MM22 VDD 7 QN VDD P l=0.18u w=1.5u 
MM21 VDD 8 7 VDD P l=0.18u w=0.57u 
MM20 2 IPM VDD VDD P l=0.18u w=1u 
MM19 VDD SDN 2 VDD P l=0.18u w=1u 
MM18 VDD E 4 VDD P l=0.18u w=0.65u 
MM17 VDD 4 3 VDD P l=0.18u w=0.65u 
MM16 16 CDN VDD VDD P l=0.18u w=0.99u 
MM15 VDD D 16 VDD P l=0.18u w=0.99u 
MM13 2 IPM 17 VSS N l=0.18u w=0.67u 
MM12 17 SDN VSS VSS N l=0.18u w=1u 
MM11 IPM 3 16 VSS N l=0.18u w=0.57u 
MM10 8 4 IPM VSS N l=0.18u w=0.84u 
MM14 VSS 2 18 VSS N l=0.18u w=0.84u 
MM9 8 CDN 18 VSS N l=0.18u w=0.84u 
MM8 6 2 VSS VSS N l=0.18u w=0.84u 
MM7 Q 6 VSS VSS N l=0.18u w=1u 
MM6 QN 7 VSS VSS N l=0.188166u w=1.014u 
MM5 VSS E 4 VSS N l=0.18u w=0.5u 
MM4 VSS 4 3 VSS N l=0.18u w=0.5u 
MM3 VSS 8 7 VSS N l=0.18u w=0.84u 
MM2 19 CDN 16 VSS N l=0.18u w=0.67u 
MM1 19 D VSS VSS N l=0.18u w=0.67u 
.ENDS labhb1

.SUBCKT labhb2 Q QN  CDN D E SDN VDD VSS
MM32 VDD 2 3 VDD P l=0.18u w=0.57u 
MM31 Q 3 VDD VDD P l=0.18u w=1.5u 
MM30 VDD 3 Q VDD P l=0.18u w=1.5u 
MM29 QN 4 VDD VDD P l=0.18u w=1.5u 
MM28 QN 4 VDD VDD P l=0.18u w=1.5u 
MM27 VDD E 6 VDD P l=0.18u w=0.65u 
MM26 VDD 6 10 VDD P l=0.18u w=0.65u 
MM24 VDD 8 4 VDD P l=0.18u w=0.57u 
MM25 VDD SDN 2 VDD P l=0.18u w=1u 
MM23 2 IPM VDD VDD P l=0.18u w=1u 
MM22 VDD 2 8 VDD P l=0.18u w=0.77u 
MM21 8 10 IPM VDD P l=0.18u w=0.67u 
MM20 16 6 IPM VDD P l=0.18u w=0.72u 
MM19 VDD CDN 8 VDD P l=0.186628u w=1.032u 
MM18 16 CDN VDD VDD P l=0.18u w=0.99u 
MM17 VDD D 16 VDD P l=0.18u w=0.99u 
MM15 17 SDN VSS VSS N l=0.18u w=1u 
MM14 2 IPM 17 VSS N l=0.18u w=0.67u 
MM13 IPM 10 16 VSS N l=0.18u w=0.57u 
MM12 8 6 IPM VSS N l=0.18u w=0.84u 
MM16 VSS 2 18 VSS N l=0.18u w=0.84u 
MM11 8 CDN 18 VSS N l=0.18u w=0.84u 
MM10 VSS 3 Q VSS N l=0.186826u w=1.002u 
MM9 Q 3 VSS VSS N l=0.186826u w=1.002u 
MM8 VSS 4 QN VSS N l=0.186826u w=1.002u 
MM7 VSS 4 QN VSS N l=0.186826u w=1.002u 
MM6 3 2 VSS VSS N l=0.18u w=0.84u 
MM5 VSS E 6 VSS N l=0.18u w=0.5u 
MM4 VSS 6 10 VSS N l=0.18u w=0.5u 
MM3 4 8 VSS VSS N l=0.18u w=0.84u 
MM2 19 CDN 16 VSS N l=0.18u w=0.67u 
MM1 19 D VSS VSS N l=0.18u w=0.67u 
.ENDS labhb2

.SUBCKT lachq1 Q  CDN D E VDD VSS
MM20 11 2 IPM VDD P l=0.18u w=1u 
MM19 12 3 IPM VDD P l=0.18u w=1.2u 
MM18 11 CDN VDD VDD P l=0.186867u w=1.066u 
MM17 11 5 VDD VDD P l=0.18u w=1.05u 
MM16 VDD IPM Q VDD P l=0.1852u w=1.5u 
MM15 VDD IPM 5 VDD P l=0.18u w=0.97u 
MM14 2 3 VDD VDD P l=0.18u w=0.71u 
MM13 3 E VDD VDD P l=0.18u w=0.71u 
MM12 VDD CDN 12 VDD P l=0.18u w=1.24u 
MM11 VDD D 12 VDD P l=0.185954u w=1.31u 
MM10 12 2 IPM VSS N l=0.18u w=0.88u 
MM9 11 3 IPM VSS N l=0.18u w=0.88u 
MM8 11 CDN 13 VSS N l=0.18u w=0.88u 
MM7 13 5 VSS VSS N l=0.18u w=0.88u 
MM6 VSS IPM Q VSS N l=0.187349u w=0.996u 
MM5 VSS IPM 5 VSS N l=0.18u w=0.48u 
MM4 12 CDN 14 VSS N l=0.18u w=1.4u 
MM3 VSS D 14 VSS N l=0.18u w=1.4u 
MM2 2 3 VSS VSS N l=0.187113u w=1.164u 
MM1 3 E VSS VSS N l=0.18u w=1.09u 
.ENDS lachq1

.SUBCKT lachq2 Q  CDN D E VDD VSS
MM22 11 2 IPM VDD P l=0.18u w=1u 
MM21 IPM 3 12 VDD P l=0.18u w=1.2u 
MM20 11 CDN VDD VDD P l=0.186867u w=1.066u 
MM19 11 5 VDD VDD P l=0.18u w=1.05u 
MM17 VDD IPM 5 VDD P l=0.18u w=0.97u 
MM18 VDD IPM Q VDD P l=0.1852u w=1.5u 
MM16 Q IPM VDD VDD P l=0.1852u w=1.5u 
MM15 2 3 VDD VDD P l=0.18u w=0.71u 
MM14 VDD E 3 VDD P l=0.18u w=0.71u 
MM13 VDD CDN 12 VDD P l=0.18u w=1.24u 
MM12 VDD D 12 VDD P l=0.185954u w=1.31u 
MM11 12 2 IPM VSS N l=0.18u w=0.88u 
MM10 11 3 IPM VSS N l=0.18u w=0.88u 
MM9 11 CDN 13 VSS N l=0.18u w=0.88u 
MM8 VSS 5 13 VSS N l=0.18u w=0.88u 
MM7 VSS IPM Q VSS N l=0.187349u w=0.996u 
MM6 VSS IPM Q VSS N l=0.187349u w=0.996u 
MM5 VSS IPM 5 VSS N l=0.18u w=0.48u 
MM4 12 CDN 14 VSS N l=0.18u w=1.4u 
MM3 VSS D 14 VSS N l=0.18u w=1.4u 
MM2 2 3 VSS VSS N l=0.187113u w=1.164u 
MM1 3 E VSS VSS N l=0.18u w=1.09u 
.ENDS lachq2

.SUBCKT laclq1 Q  CDN D EN VDD VSS
MM20 IPM 2 12 VDD P l=0.18u w=0.75u 
MM19 11 3 IPM VDD P l=0.18u w=0.75u 
MM18 11 CDN VDD VDD P l=0.186564u w=1.042u 
MM17 11 5 VDD VDD P l=0.18729u w=1.07u 
MM16 VDD IPM 5 VDD P l=0.18u w=0.52u 
MM15 VDD IPM Q VDD P l=0.18u w=1.54u 
MM14 VDD 3 2 VDD P l=0.18u w=0.68u 
MM13 VDD EN 3 VDD P l=0.18u w=0.68u 
MM12 VDD CDN 12 VDD P l=0.18u w=1.14u 
MM11 VDD D 12 VDD P l=0.188862u w=1.239u 
MM10 IPM 2 11 VSS N l=0.18u w=0.6u 
MM9 IPM 3 12 VSS N l=0.18u w=0.6u 
MM8 13 CDN 11 VSS N l=0.18u w=0.75u 
MM7 VSS 5 13 VSS N l=0.18u w=0.75u 
MM6 VSS IPM 5 VSS N l=0.18u w=0.48u 
MM5 VSS IPM Q VSS N l=0.18u w=1.04u 
MM4 14 CDN 12 VSS N l=0.18u w=0.77u 
MM3 14 D VSS VSS N l=0.18u w=0.77u 
MM2 VSS 3 2 VSS N l=0.18u w=0.52u 
MM1 3 EN VSS VSS N l=0.18u w=0.52u 
.ENDS laclq1

.SUBCKT laclq2 Q  CDN D EN VDD VSS
MM22 6 2 12 VDD P l=0.18u w=1.01u 
MM21 11 CDN VDD VDD P l=0.18828u w=1.058u 
MM20 6 4 11 VDD P l=0.18u w=1.01u 
MM19 11 5 VDD VDD P l=0.18u w=1u 
MM18 VDD 6 5 VDD P l=0.18u w=0.61u 
MM17 VDD 6 Q VDD P l=0.18u w=1.5u 
MM16 Q 6 VDD VDD P l=0.18u w=1.5u 
MM15 VDD 4 2 VDD P l=0.18u w=0.55u 
MM14 VDD EN 4 VDD P l=0.18u w=0.65u 
MM13 12 CDN VDD VDD P l=0.18u w=1.03u 
MM12 12 D VDD VDD P l=0.1875u w=1.104u 
MM11 6 2 11 VSS N l=0.18u w=0.81u 
MM10 13 CDN 11 VSS N l=0.18u w=0.72u 
MM9 12 4 6 VSS N l=0.18u w=0.81u 
MM8 13 5 VSS VSS N l=0.18u w=0.72u 
MM7 VSS 6 5 VSS N l=0.18u w=0.84u 
MM6 VSS 6 Q VSS N l=0.18u w=1u 
MM5 VSS 6 Q VSS N l=0.18u w=1u 
MM4 VSS 4 2 VSS N l=0.18u w=0.5u 
MM3 4 EN VSS VSS N l=0.18u w=0.5u 
MM2 14 CDN 12 VSS N l=0.18u w=0.74u 
MM1 VSS D 14 VSS N l=0.18u w=0.74u 
.ENDS laclq2

.SUBCKT lanhb1 Q QN  D E VDD VSS
MM18 4 E VDD VDD P l=0.18u w=0.84u 
MM17 10 3 IPM VDD P l=0.18u w=0.5u 
MM15 12 4 IPM VDD P l=0.1865u w=1.2u 
MM16 VDD 4 3 VDD P l=0.18806u w=1.206u 
MM12 VDD D 12 VDD P l=0.192908u w=1.269u 
MM14 VDD IPM 6 VDD P l=0.18u w=1.54u 
MM13 VDD 6 10 VDD P l=0.18u w=0.5u 
MM11 Q IPM VDD VDD P l=0.18u w=1.5u 
MM10 QN 6 VDD VDD P l=0.18u w=1.5u 
MM9 IPM 3 12 VSS N l=0.185787u w=1.182u 
MM7 IPM 4 10 VSS N l=0.18u w=0.8u 
MM8 3 4 VSS VSS N l=0.185787u w=1.182u 
MM6 6 IPM VSS VSS N l=0.18u w=0.84u 
MM5 VSS 6 10 VSS N l=0.18u w=0.8u 
MM4 VSS D 12 VSS N l=0.186172u w=1.186u 
MM3 VSS IPM Q VSS N l=0.186826u w=1.002u 
MM2 VSS 6 QN VSS N l=0.186826u w=1.002u 
MM1 4 E VSS VSS N l=0.18u w=0.53u 
.ENDS lanhb1

.SUBCKT lanhb2 Q QN  D E VDD VSS
MM22 7 E VDD VDD P l=0.18u w=0.84u 
MM19 IPM 5 11 VDD P l=0.18u w=0.5u 
MM16 12 7 IPM VDD P l=0.18u w=1.2u 
MM20 VDD IPM 3 VDD P l=0.18u w=1.54u 
MM21 VDD 3 11 VDD P l=0.18u w=0.5u 
MM17 VDD 7 5 VDD P l=0.185691u w=1.202u 
MM18 VDD D 12 VDD P l=0.18922u w=1.243u 
MM15 QN 3 VDD VDD P l=0.18u w=1.5u 
MM14 VDD 3 QN VDD P l=0.18u w=1.5u 
MM13 Q IPM VDD VDD P l=0.18u w=1.5u 
MM12 VDD IPM Q VDD P l=0.18u w=1.5u 
MM10 3 IPM VSS VSS N l=0.18u w=0.84u 
MM9 VSS D 12 VSS N l=0.185787u w=1.182u 
MM8 IPM 5 12 VSS N l=0.185787u w=1.182u 
MM6 IPM 7 11 VSS N l=0.18u w=0.8u 
MM7 5 7 VSS VSS N l=0.185787u w=1.182u 
MM11 11 3 VSS VSS N l=0.18u w=0.8u 
MM5 VSS 3 QN VSS N l=0.186826u w=1.002u 
MM4 VSS 3 QN VSS N l=0.186826u w=1.002u 
MM3 VSS IPM Q VSS N l=0.186826u w=1.002u 
MM2 VSS IPM Q VSS N l=0.186826u w=1.002u 
MM1 7 E VSS VSS N l=0.18u w=0.53u 
.ENDS lanhb2

.SUBCKT lanhn1 QN  D E VDD VSS
MM18 12 2 IPM VDD P l=0.18u w=0.65u 
MM17 IPM 3 9 VDD P l=0.18u w=0.7u 
MM16 12 4 VDD VDD P l=0.18u w=0.65u 
MM15 4 IPM VDD VDD P l=0.18u w=0.6u 
MM14 VDD 6 9 VDD P l=0.18u w=0.7u 
MM13 QN IPM VDD VDD P l=0.18u w=1.5u 
MM12 3 E VDD VDD P l=0.18u w=0.52u 
MM11 VDD 3 2 VDD P l=0.18u w=0.52u 
MM10 VDD D 6 VDD P l=0.18u w=0.52u 
MM8 12 3 IPM VSS N l=0.18u w=0.57u 
MM7 12 4 VSS VSS N l=0.18u w=0.57u 
MM9 9 2 IPM VSS N l=0.18u w=0.57u 
MM6 4 IPM VSS VSS N l=0.18u w=0.57u 
MM5 9 6 VSS VSS N l=0.18u w=0.57u 
MM4 QN IPM VSS VSS N l=0.18u w=1u 
MM3 3 E VSS VSS N l=0.18u w=0.48u 
MM2 VSS 3 2 VSS N l=0.18u w=0.48u 
MM1 VSS D 6 VSS N l=0.18u w=0.48u 
.ENDS lanhn1

.SUBCKT lanhn2 QN  D E VDD VSS
MM20 11 2 IPM VDD P l=0.18u w=0.65u 
MM19 IPM 3 12 VDD P l=0.18u w=0.7u 
MM18 11 4 VDD VDD P l=0.18u w=0.65u 
MM17 4 IPM VDD VDD P l=0.18u w=0.6u 
MM16 VDD 6 12 VDD P l=0.18u w=0.7u 
MM15 QN IPM VDD VDD P l=0.18u w=1.5u 
MM14 QN IPM VDD VDD P l=0.18u w=1.5u 
MM13 3 E VDD VDD P l=0.18u w=0.52u 
MM12 VDD 3 2 VDD P l=0.18u w=0.52u 
MM11 VDD D 6 VDD P l=0.18u w=0.52u 
MM9 11 3 IPM VSS N l=0.18u w=0.57u 
MM8 VSS 4 11 VSS N l=0.18u w=0.57u 
MM10 12 2 IPM VSS N l=0.18u w=0.57u 
MM7 VSS IPM 4 VSS N l=0.18u w=0.57u 
MM6 12 6 VSS VSS N l=0.18u w=0.57u 
MM5 QN IPM VSS VSS N l=0.18u w=1u 
MM4 QN IPM VSS VSS N l=0.18u w=1u 
MM3 3 E VSS VSS N l=0.18u w=0.48u 
MM2 VSS 3 2 VSS N l=0.18u w=0.48u 
MM1 VSS D 6 VSS N l=0.18u w=0.48u 
.ENDS lanhn2

.SUBCKT lanhq1 Q  D E VDD VSS
MM16 4 E VDD VDD P l=0.18u w=0.68u 
MM15 10 3 IPM VDD P l=0.18u w=0.6u 
MM12 10 5 VDD VDD P l=0.18u w=0.52u 
MM14 11 4 IPM VDD P l=0.18u w=0.82u 
MM13 VDD 4 3 VDD P l=0.18u w=0.68u 
MM11 VDD IPM 5 VDD P l=0.18u w=0.52u 
MM10 VDD D 11 VDD P l=0.18u w=0.82u 
MM9 Q IPM VDD VDD P l=0.18u w=1.51u 
MM7 VSS 4 3 VSS N l=0.18u w=0.54u 
MM8 IPM 3 11 VSS N l=0.18u w=0.88u 
MM6 10 4 IPM VSS N l=0.18u w=0.88u 
MM5 10 5 VSS VSS N l=0.18u w=0.88u 
MM4 5 IPM VSS VSS N l=0.18u w=0.88u 
MM3 VSS D 11 VSS N l=0.18u w=0.88u 
MM2 VSS IPM Q VSS N l=0.18u w=1u 
MM1 4 E VSS VSS N l=0.18u w=0.5u 
.ENDS lanhq1

.SUBCKT lanhq2 Q  D E VDD VSS
MM18 6 E VDD VDD P l=0.18u w=0.68u 
MM17 10 3 IPM VDD P l=0.18u w=0.6u 
MM16 10 4 VDD VDD P l=0.18u w=0.52u 
MM15 VDD IPM 4 VDD P l=0.18u w=0.52u 
MM14 11 6 IPM VDD P l=0.18u w=0.82u 
MM13 VDD 6 3 VDD P l=0.18u w=0.68u 
MM12 VDD D 11 VDD P l=0.18u w=0.82u 
MM11 Q IPM VDD VDD P l=0.184554u w=1.502u 
MM10 VDD IPM Q VDD P l=0.184861u w=1.506u 
MM7 4 IPM VSS VSS N l=0.18u w=0.88u 
MM6 VSS 6 3 VSS N l=0.18u w=0.54u 
MM8 10 4 VSS VSS N l=0.18u w=0.88u 
MM5 10 6 IPM VSS N l=0.18u w=0.88u 
MM9 IPM 3 11 VSS N l=0.18u w=0.88u 
MM4 VSS D 11 VSS N l=0.18u w=0.88u 
MM3 VSS IPM Q VSS N l=0.187276u w=1.006u 
MM2 VSS IPM Q VSS N l=0.186826u w=1.002u 
MM1 6 E VSS VSS N l=0.18u w=0.5u 
.ENDS lanhq2

.SUBCKT lanht1 Z  D E OE VDD VSS
MM20 VDD 2 6 VDD P l=0.18u w=0.68u 
MM19 13 2 nint VDD P l=0.18u w=0.82u 
MM15 12 6 nint VDD P l=0.18u w=0.6u 
MM17 VDD nint 3 VDD P l=0.18u w=0.52u 
MM16 13 D VDD VDD P l=0.18u w=0.82u 
MM18 VDD 3 12 VDD P l=0.18u w=0.52u 
MM14 8 OE VDD VDD P l=0.18u w=0.82u 
MM12 15 nint Z VDD P l=0.18u w=1.5u 
MM13 15 8 VDD VDD P l=0.18u w=1.5u 
MM11 2 E VDD VDD P l=0.18u w=0.68u 
MM10 VSS 2 6 VSS N l=0.18u w=0.54u 
MM9 12 2 nint VSS N l=0.18u w=0.44u 
MM8 12 3 VSS VSS N l=0.18u w=0.44u 
MM7 3 nint VSS VSS N l=0.18u w=0.44u 
MM5 nint 6 13 VSS N l=0.18u w=0.6u 
MM6 VSS D 13 VSS N l=0.18u w=0.6u 
MM4 8 OE VSS VSS N l=0.18u w=0.63u 
MM2 Z nint 14 VSS N l=0.18u w=1u 
MM3 14 OE VSS VSS N l=0.18u w=1u 
MM1 VSS E 2 VSS N l=0.18u w=0.5u 
.ENDS lanht1

.SUBCKT lanht2 Z  D E OE VDD VSS
MM21 VDD 5 6 VDD P l=0.18u w=0.68u 
MM24 VDD nint 3 VDD P l=0.18u w=0.52u 
MM20 13 5 nint VDD P l=0.18u w=0.82u 
MM19 12 6 nint VDD P l=0.18u w=0.6u 
MM22 13 D VDD VDD P l=0.18u w=0.82u 
MM23 VDD 3 12 VDD P l=0.18u w=0.52u 
MM18 VDD nint 16 VDD P l=0.18u w=1.5u 
MM17 Z 7 16 VDD P l=0.18u w=1.5u 
MM15 7 OE VDD VDD P l=0.186341u w=1.23u 
MM14 17 7 Z VDD P l=0.18u w=1.5u 
MM16 17 nint VDD VDD P l=0.18u w=1.5u 
MM13 5 E VDD VDD P l=0.18u w=0.68u 
MM12 VSS nint 3 VSS N l=0.18u w=0.44u 
MM11 VSS 3 12 VSS N l=0.18u w=0.44u 
MM9 12 5 nint VSS N l=0.18u w=0.44u 
MM8 VSS 5 6 VSS N l=0.18u w=0.54u 
MM7 nint 6 13 VSS N l=0.18u w=0.6u 
MM10 VSS D 13 VSS N l=0.18u w=0.6u 
MM5 Z OE 14 VSS N l=0.18u w=1u 
MM6 VSS nint 14 VSS N l=0.18u w=1u 
MM4 VSS E 5 VSS N l=0.18u w=0.5u 
MM2 VSS OE 7 VSS N l=0.18u w=0.94u 
MM1 15 OE Z VSS N l=0.18u w=1u 
MM3 15 nint VSS VSS N l=0.18u w=1u 
.ENDS lanht2

.SUBCKT lanlb1 Q QN  D EN VDD VSS
MM18 4 EN VDD VDD P l=0.18u w=0.57u 
MM17 12 3 IPM VDD P l=0.18u w=0.72u 
MM16 11 4 IPM VDD P l=0.18u w=0.6u 
MM15 3 4 VDD VDD P l=0.18u w=1.12u 
MM14 VDD 5 11 VDD P l=0.18u w=0.72u 
MM13 VDD IPM 5 VDD P l=0.18u w=0.72u 
MM12 VDD D 12 VDD P l=0.18u w=0.93u 
MM11 QN 5 VDD VDD P l=0.184554u w=1.502u 
MM10 Q IPM VDD VDD P l=0.184554u w=1.502u 
MM8 3 4 VSS VSS N l=0.18u w=0.58u 
MM9 IPM 3 11 VSS N l=0.18u w=0.55u 
MM7 IPM 4 12 VSS N l=0.18u w=0.55u 
MM6 VSS 5 11 VSS N l=0.18u w=0.55u 
MM5 5 IPM VSS VSS N l=0.18u w=0.67u 
MM4 VSS D 12 VSS N l=0.18u w=0.94u 
MM2 Q IPM VSS VSS N l=0.186826u w=1.002u 
MM3 QN 5 VSS VSS N l=0.186826u w=1.002u 
MM1 4 EN VSS VSS N l=0.18u w=0.84u 
.ENDS lanlb1

.SUBCKT lanlb2 Q QN  D EN VDD VSS
MM22 6 EN VDD VDD P l=0.18u w=0.57u 
MM21 VDD 3 11 VDD P l=0.18u w=0.72u 
MM18 11 6 IPM VDD P l=0.18u w=0.6u 
MM20 VDD IPM 3 VDD P l=0.18u w=0.72u 
MM19 12 5 IPM VDD P l=0.18u w=0.72u 
MM17 VDD 6 5 VDD P l=0.18u w=1.12u 
MM16 VDD D 12 VDD P l=0.18u w=0.93u 
MM15 VDD 3 QN VDD P l=0.184554u w=1.502u 
MM14 QN 3 VDD VDD P l=0.184554u w=1.502u 
MM13 VDD IPM Q VDD P l=0.184554u w=1.502u 
MM12 VDD IPM Q VDD P l=0.184554u w=1.502u 
MM10 3 IPM VSS VSS N l=0.18u w=0.67u 
MM9 VSS D 12 VSS N l=0.18u w=0.94u 
MM6 IPM 6 12 VSS N l=0.18u w=0.55u 
MM11 VSS 3 11 VSS N l=0.18u w=0.55u 
MM8 IPM 5 11 VSS N l=0.18u w=0.55u 
MM7 5 6 VSS VSS N l=0.18u w=0.58u 
MM5 VSS 3 QN VSS N l=0.186826u w=1.002u 
MM4 VSS 3 QN VSS N l=0.186826u w=1.002u 
MM3 VSS IPM Q VSS N l=0.186826u w=1.002u 
MM2 VSS IPM Q VSS N l=0.186826u w=1.002u 
MM1 6 EN VSS VSS N l=0.18u w=0.84u 
.ENDS lanlb2

.SUBCKT lanln1 QN  D EN VDD VSS
MM18 IPM 2 9 VDD P l=0.18u w=1.03u 
MM17 IPM 3 12 VDD P l=0.18u w=0.6u 
MM16 VDD 4 12 VDD P l=0.18u w=0.52u 
MM15 VDD IPM 4 VDD P l=0.18u w=0.52u 
MM14 9 6 VDD VDD P l=0.189333u w=1.125u 
MM13 QN IPM VDD VDD P l=0.18u w=1.5u 
MM12 VDD EN 3 VDD P l=0.18u w=0.68u 
MM11 2 3 VDD VDD P l=0.18u w=0.68u 
MM10 6 D VDD VDD P l=0.18u w=0.52u 
MM9 IPM 2 12 VSS N l=0.18u w=0.57u 
MM7 12 4 VSS VSS N l=0.18u w=0.48u 
MM8 9 3 IPM VSS N l=0.18u w=0.72u 
MM5 9 6 VSS VSS N l=0.18u w=0.75u 
MM6 4 IPM VSS VSS N l=0.18u w=0.48u 
MM4 QN IPM VSS VSS N l=0.18u w=1u 
MM3 VSS EN 3 VSS N l=0.18u w=0.52u 
MM2 VSS 3 2 VSS N l=0.18u w=0.52u 
MM1 VSS D 6 VSS N l=0.18u w=0.48u 
.ENDS lanln1

.SUBCKT lanln2 QN  D EN VDD VSS
MM20 IPM 2 12 VDD P l=0.18u w=1.03u 
MM19 IPM 3 11 VDD P l=0.18u w=0.6u 
MM18 VDD 4 11 VDD P l=0.18u w=0.52u 
MM17 VDD IPM 4 VDD P l=0.18u w=0.52u 
MM16 12 6 VDD VDD P l=0.189333u w=1.125u 
MM15 VDD IPM QN VDD P l=0.185469u w=1.514u 
MM14 QN IPM VDD VDD P l=0.18u w=1.44u 
MM13 VDD EN 3 VDD P l=0.18u w=0.68u 
MM12 2 3 VDD VDD P l=0.18u w=0.68u 
MM11 6 D VDD VDD P l=0.18u w=0.52u 
MM10 IPM 2 11 VSS N l=0.18u w=0.57u 
MM8 VSS 4 11 VSS N l=0.18u w=0.48u 
MM9 12 3 IPM VSS N l=0.18u w=0.72u 
MM6 12 6 VSS VSS N l=0.18u w=0.75u 
MM7 VSS IPM 4 VSS N l=0.18u w=0.48u 
MM5 VSS IPM QN VSS N l=0.187276u w=1.006u 
MM4 QN IPM VSS VSS N l=0.18u w=1u 
MM3 VSS EN 3 VSS N l=0.18u w=0.52u 
MM2 VSS 3 2 VSS N l=0.18u w=0.52u 
MM1 VSS D 6 VSS N l=0.18u w=0.48u 
.ENDS lanln2

.SUBCKT lanlq1 Q  D EN VDD VSS
MM16 4 EN VDD VDD P l=0.18u w=0.6u 
MM14 3 4 VDD VDD P l=0.18u w=0.68u 
MM13 10 4 IPM VDD P l=0.18u w=0.78u 
MM12 10 5 VDD VDD P l=0.18u w=0.52u 
MM15 IPM 3 11 VDD P l=0.18u w=0.78u 
MM11 5 IPM VDD VDD P l=0.18u w=0.52u 
MM10 11 D VDD VDD P l=0.186042u w=1.132u 
MM9 Q IPM VDD VDD P l=0.18u w=1.5u 
MM7 VSS 4 3 VSS N l=0.18u w=0.84u 
MM8 IPM 3 10 VSS N l=0.18u w=0.6u 
MM6 11 4 IPM VSS N l=0.18u w=0.6u 
MM5 VSS 5 10 VSS N l=0.18u w=0.79u 
MM4 VSS IPM 5 VSS N l=0.18u w=0.79u 
MM3 VSS D 11 VSS N l=0.187205u w=1.016u 
MM2 VSS IPM Q VSS N l=0.18u w=1u 
MM1 4 EN VSS VSS N l=0.18u w=0.48u 
.ENDS lanlq1

.SUBCKT lanlq2 Q  D EN VDD VSS
MM18 6 EN VDD VDD P l=0.18u w=0.6u 
MM16 3 IPM VDD VDD P l=0.18u w=0.52u 
MM14 5 6 VDD VDD P l=0.18u w=0.68u 
MM17 10 3 VDD VDD P l=0.18u w=0.52u 
MM13 10 6 IPM VDD P l=0.18u w=0.78u 
MM15 IPM 5 11 VDD P l=0.18u w=0.78u 
MM12 11 D VDD VDD P l=0.186042u w=1.132u 
MM11 Q IPM VDD VDD P l=0.185469u w=1.514u 
MM10 Q IPM VDD VDD P l=0.18u w=1.44u 
MM9 VSS 3 10 VSS N l=0.18u w=0.79u 
MM6 IPM 5 10 VSS N l=0.18u w=0.6u 
MM8 VSS IPM 3 VSS N l=0.18u w=0.79u 
MM5 VSS 6 5 VSS N l=0.18u w=0.84u 
MM7 VSS D 11 VSS N l=0.187205u w=1.016u 
MM4 11 6 IPM VSS N l=0.18u w=0.6u 
MM3 VSS IPM Q VSS N l=0.187276u w=1.006u 
MM2 VSS IPM Q VSS N l=0.18u w=1u 
MM1 6 EN VSS VSS N l=0.18u w=0.48u 
.ENDS lanlq2

.SUBCKT mffnrb1 Q QN  CP D ENN VDD VSS
MM36 20 2 5 VDD P l=0.18u w=0.6u 
MM35 17 3 5 VDD P l=0.18u w=0.6u 
MM34 17 4 VDD VDD P l=0.18u w=0.71u 
MM33 VDD 5 4 VDD P l=0.18u w=1.35u 
MM32 6 2 8 VDD P l=0.18u w=0.65u 
MM29 VDD 7 8 VDD P l=0.18u w=0.52u 
MM31 4 3 6 VDD P l=0.18854u w=1.082u 
MM30 VDD 6 7 VDD P l=0.18671u w=1.234u 
MM28 19 8 VDD VDD P l=0.18u w=0.5u 
MM23 19 12 20 VDD P l=0.18u w=0.6u 
MM27 VDD CP 3 VDD P l=0.18u w=0.68u 
MM26 VDD 3 2 VDD P l=0.18u w=0.68u 
MM25 VDD D 18 VDD P l=0.18u w=0.52u 
MM24 18 11 20 VDD P l=0.18u w=0.6u 
MM22 VDD 12 11 VDD P l=0.18u w=0.52u 
MM21 VDD ENN 12 VDD P l=0.18u w=0.52u 
MM20 VDD 6 QN VDD P l=0.18u w=1.5u 
MM19 VDD 7 Q VDD P l=0.18u w=1.5u 
MM18 17 2 5 VSS N l=0.18u w=0.65u 
MM16 VSS 4 17 VSS N l=0.18u w=0.37u 
MM17 6 2 4 VSS N l=0.18u w=1.26u 
MM15 8 3 6 VSS N l=0.18u w=0.84u 
MM13 8 7 VSS VSS N l=0.18u w=0.51u 
MM14 VSS 5 4 VSS N l=0.186207u w=1.334u 
MM12 5 3 20 VSS N l=0.18u w=0.65u 
MM11 7 6 VSS VSS N l=0.189002u w=1.273u 
MM10 VSS ENN 12 VSS N l=0.18u w=0.43u 
MM9 19 8 VSS VSS N l=0.18u w=0.43u 
MM5 19 11 20 VSS N l=0.18u w=0.84u 
MM8 VSS CP 3 VSS N l=0.18u w=0.6u 
MM7 VSS 3 2 VSS N l=0.18u w=0.51u 
MM4 VSS 12 11 VSS N l=0.18u w=0.49u 
MM3 18 12 20 VSS N l=0.18u w=0.84u 
MM6 18 D VSS VSS N l=0.18u w=0.84u 
MM2 QN 6 VSS VSS N l=0.18u w=1u 
MM1 Q 7 VSS VSS N l=0.18u w=1u 
.ENDS mffnrb1

.SUBCKT mffnrb2 Q QN  CP D ENN VDD VSS
MM40 20 2 4 VDD P l=0.18u w=0.6u 
MM39 17 3 VDD VDD P l=0.18u w=0.71u 
MM37 17 5 4 VDD P l=0.18u w=0.6u 
MM38 VDD 4 3 VDD P l=0.18u w=1.35u 
MM36 6 2 8 VDD P l=0.18u w=0.65u 
MM30 VDD 7 8 VDD P l=0.18u w=0.52u 
MM32 3 5 6 VDD P l=0.18854u w=1.082u 
MM35 VDD 6 QN VDD P l=0.184554u w=1.502u 
MM34 VDD 6 QN VDD P l=0.184861u w=1.506u 
MM33 VDD 6 7 VDD P l=0.185971u w=1.226u 
MM31 VDD 7 Q VDD P l=0.184554u w=1.502u 
MM29 VDD 7 Q VDD P l=0.184861u w=1.506u 
MM28 19 8 VDD VDD P l=0.18u w=0.5u 
MM23 19 12 20 VDD P l=0.18u w=0.6u 
MM27 VDD CP 5 VDD P l=0.18u w=0.68u 
MM26 VDD 5 2 VDD P l=0.18u w=0.68u 
MM25 VDD D 18 VDD P l=0.18u w=0.52u 
MM24 18 11 20 VDD P l=0.18u w=0.6u 
MM22 VDD 12 11 VDD P l=0.18u w=0.52u 
MM21 VDD ENN 12 VDD P l=0.18u w=0.52u 
MM20 17 2 4 VSS N l=0.18u w=0.65u 
MM18 VSS 3 17 VSS N l=0.18u w=0.37u 
MM19 6 2 3 VSS N l=0.18u w=1.26u 
MM17 8 5 6 VSS N l=0.18u w=0.84u 
MM15 VSS 7 8 VSS N l=0.18u w=0.51u 
MM16 VSS 4 3 VSS N l=0.186207u w=1.334u 
MM14 4 5 20 VSS N l=0.18u w=0.65u 
MM13 VSS 6 QN VSS N l=0.187276u w=1.006u 
MM12 QN 6 VSS VSS N l=0.186826u w=1.002u 
MM11 VSS 6 7 VSS N l=0.18u w=1.27u 
MM10 VSS 7 Q VSS N l=0.187276u w=1.006u 
MM9 VSS 7 Q VSS N l=0.186826u w=1.002u 
MM8 VSS ENN 12 VSS N l=0.18u w=0.43u 
MM7 19 8 VSS VSS N l=0.18u w=0.43u 
MM3 19 11 20 VSS N l=0.18u w=0.84u 
MM6 VSS CP 5 VSS N l=0.18u w=0.6u 
MM5 VSS 5 2 VSS N l=0.18u w=0.51u 
MM2 VSS 12 11 VSS N l=0.18u w=0.49u 
MM1 18 12 20 VSS N l=0.18u w=0.84u 
MM4 18 D VSS VSS N l=0.18u w=0.84u 
.ENDS mffnrb2

.SUBCKT mi02d0 S ZN  I0 I1 VDD VSS
MM14 7 2 VDD VDD P l=0.18u w=0.79u 
MM12 12 4 2 VDD P l=0.188782u w=1.141u 
MM10 2 S 13 VDD P l=0.18u w=0.79u 
MM11 12 I1 VDD VDD P l=0.18u w=1.05u 
MM13 VDD I0 13 VDD P l=0.18u w=0.79u 
MM9 VDD S 4 VDD P l=0.18u w=0.54u 
MM8 ZN 7 VDD VDD P l=0.18u w=0.73u 
MM5 VSS 7 ZN VSS N l=0.18u w=0.42u 
MM7 7 2 VSS VSS N l=0.18u w=0.42u 
MM6 VSS I0 10 VSS N l=0.18u w=0.98u 
MM4 2 4 10 VSS N l=0.18u w=0.98u 
MM2 VSS S 4 VSS N l=0.18u w=0.48u 
MM1 2 S 11 VSS N l=0.18u w=0.98u 
MM3 11 I1 VSS VSS N l=0.18u w=0.98u 
.ENDS mi02d0

.SUBCKT mi02d1 S ZN  I0 I1 VDD VSS
MM14 VDD 2 7 VDD P l=0.18u w=0.79u 
MM12 12 4 2 VDD P l=0.188127u w=1.196u 
MM9 13 S 2 VDD P l=0.18u w=0.79u 
MM11 12 I1 VDD VDD P l=0.18u w=1.11u 
MM10 4 S VDD VDD P l=0.18661u w=1.18u 
MM13 13 I0 VDD VDD P l=0.18u w=0.79u 
MM8 ZN 7 VDD VDD P l=0.184968u w=1.57u 
MM7 7 2 VSS VSS N l=0.18u w=0.42u 
MM6 VSS I0 10 VSS N l=0.18u w=0.98u 
MM5 2 4 10 VSS N l=0.18u w=0.98u 
MM3 4 S VSS VSS N l=0.18661u w=1.18u 
MM2 2 S 11 VSS N l=0.18u w=1.11u 
MM4 11 I1 VSS VSS N l=0.18u w=1.11u 
MM1 VSS 7 ZN VSS N l=0.18661u w=1.18u 
.ENDS mi02d1

.SUBCKT mi02d2 S ZN  I0 I1 VDD VSS
MM15 VDD 3 7 VDD P l=0.18u w=0.79u 
MM14 12 4 3 VDD P l=0.188127u w=1.196u 
MM11 13 S 3 VDD P l=0.18u w=0.79u 
MM13 12 I1 VDD VDD P l=0.18u w=1.11u 
MM12 4 S VDD VDD P l=0.18661u w=1.18u 
MM16 VDD I0 13 VDD P l=0.18u w=0.79u 
MM10 ZN 7 VDD VDD P l=0.185098u w=1.53u 
MM9 ZN 7 VDD VDD P l=0.18u w=1.46u 
MM7 7 3 VSS VSS N l=0.18u w=0.42u 
MM8 VSS I0 10 VSS N l=0.18u w=0.98u 
MM6 3 4 10 VSS N l=0.18u w=0.98u 
MM4 4 S VSS VSS N l=0.18661u w=1.18u 
MM3 3 S 11 VSS N l=0.18u w=1.11u 
MM5 11 I1 VSS VSS N l=0.18u w=1.11u 
MM2 VSS 7 ZN VSS N l=0.18661u w=1.18u 
MM1 VSS 7 ZN VSS N l=0.18u w=1.11u 
.ENDS mi02d2

.SUBCKT mi02d4 S ZN  I0 I1 VDD VSS
MM18 VDD 2 7 VDD P l=0.18u w=0.79u 
MM16 12 4 2 VDD P l=0.188127u w=1.196u 
MM13 13 S 2 VDD P l=0.18u w=0.79u 
MM15 12 I1 VDD VDD P l=0.18u w=1.11u 
MM14 4 S VDD VDD P l=0.18661u w=1.18u 
MM17 13 I0 VDD VDD P l=0.18u w=0.79u 
MM12 ZN 7 VDD VDD P l=0.183786u w=2.06u 
MM11 ZN 7 VDD VDD P l=0.18u w=1.99u 
MM10 ZN 7 VDD VDD P l=0.18u w=1.99u 
MM9 7 2 VSS VSS N l=0.18u w=0.42u 
MM8 VSS I0 10 VSS N l=0.18u w=0.98u 
MM7 2 4 10 VSS N l=0.18u w=0.98u 
MM5 4 S VSS VSS N l=0.18661u w=1.18u 
MM4 2 S 11 VSS N l=0.18u w=1.11u 
MM6 11 I1 VSS VSS N l=0.18u w=1.11u 
MM3 ZN 7 VSS VSS N l=0.184643u w=1.68u 
MM2 ZN 7 VSS VSS N l=0.18u w=1.61u 
MM1 VSS 7 ZN VSS N l=0.18u w=1.61u 
.ENDS mi02d4

.SUBCKT mx02d0 S Z  I0 I1 VDD VSS
MM12 12 2 5 VDD P l=0.18u w=0.77u 
MM10 11 S 5 VDD P l=0.18u w=0.68u 
MM11 2 S VDD VDD P l=0.18u w=0.52u 
MM9 VDD I0 11 VDD P l=0.18u w=0.68u 
MM8 VDD 5 Z VDD P l=0.18u w=0.93u 
MM7 12 I1 VDD VDD P l=0.18u w=0.77u 
MM5 VSS S 2 VSS N l=0.18u w=0.48u 
MM6 9 2 5 VSS N l=0.18u w=0.88u 
MM4 10 S 5 VSS N l=0.18u w=0.88u 
MM3 9 I0 VSS VSS N l=0.18u w=0.88u 
MM2 Z 5 VSS VSS N l=0.18u w=0.88u 
MM1 10 I1 VSS VSS N l=0.18u w=0.88u 
.ENDS mx02d0

.SUBCKT mx02d1 S Z  I0 I1 VDD VSS
MM12 12 2 4 VDD P l=0.18u w=1.34u 
MM11 11 S 4 VDD P l=0.186178u w=1.418u 
MM10 2 S VDD VDD P l=0.18u w=0.63u 
MM9 VDD 4 Z VDD P l=0.18u w=1.34u 
MM8 11 I0 VDD VDD P l=0.185532u w=1.41u 
MM7 12 I1 VDD VDD P l=0.18u w=1.34u 
MM5 2 S VSS VSS N l=0.18u w=0.55u 
MM6 9 2 4 VSS N l=0.187027u w=1.11u 
MM4 10 S 4 VSS N l=0.18u w=1.04u 
MM3 Z 4 VSS VSS N l=0.187027u w=1.11u 
MM2 9 I0 VSS VSS N l=0.18u w=1.04u 
MM1 VSS I1 10 VSS N l=0.18u w=1.04u 
.ENDS mx02d1

.SUBCKT mx02d2 S Z  I0 I1 VDD VSS
MM14 12 2 4 VDD P l=0.18u w=1.4u 
MM13 11 S 4 VDD P l=0.185617u w=1.474u 
MM12 VDD S 2 VDD P l=0.18u w=0.63u 
MM11 VDD 4 Z VDD P l=0.185306u w=1.47u 
MM10 VDD 4 Z VDD P l=0.18u w=1.4u 
MM9 11 I0 VDD VDD P l=0.185306u w=1.47u 
MM8 12 I1 VDD VDD P l=0.18u w=1.4u 
MM6 2 S VSS VSS N l=0.18u w=0.55u 
MM7 9 2 4 VSS N l=0.187433u w=1.114u 
MM5 10 S 4 VSS N l=0.18u w=1.04u 
MM4 Z 4 VSS VSS N l=0.186935u w=1.194u 
MM3 Z 4 VSS VSS N l=0.18u w=1.12u 
MM2 VSS I0 9 VSS N l=0.18u w=1.12u 
MM1 VSS I1 10 VSS N l=0.18u w=1.04u 
.ENDS mx02d2

.SUBCKT mx02d4 S Z  I0 I1 VDD VSS
MM15 VDD 3 Z VDD P l=0.185306u w=1.47u 
MM14 VDD 3 Z VDD P l=0.18u w=1.4u 
MM13 VDD 3 Z VDD P l=0.18u w=1.4u 
MM12 11 4 3 VDD P l=0.18u w=1.4u 
MM11 11 I1 VDD VDD P l=0.18u w=1.4u 
MM10 12 S 3 VDD P l=0.185617u w=1.474u 
MM16 12 I0 VDD VDD P l=0.185306u w=1.47u 
MM9 VDD S 4 VDD P l=0.18u w=0.63u 
MM6 Z 3 VSS VSS N l=0.186935u w=1.194u 
MM7 Z 3 VSS VSS N l=0.186935u w=1.194u 
MM5 Z 3 VSS VSS N l=0.18u w=1.12u 
MM4 9 4 3 VSS N l=0.186172u w=1.186u 
MM1 10 S 3 VSS N l=0.18u w=1.04u 
MM8 VSS I0 9 VSS N l=0.18u w=1.12u 
MM2 VSS S 4 VSS N l=0.18u w=0.55u 
MM3 10 I1 VSS VSS N l=0.18u w=1.04u 
.ENDS mx02d4

.SUBCKT mx04d0 Z  I0 I1 I2 I3 S0 S1 VDD VSS
MM30 21 I2 VDD VDD P l=0.18u w=1.06u 
MM29 27 3 21 VDD P l=0.18u w=1.06u 
MM25 VDD 5 Z VDD P l=0.18u w=0.68u 
MM28 22 3 24 VDD P l=0.18u w=1.06u 
MM24 22 I3 VDD VDD P l=0.18u w=1.06u 
MM26 23 S1 25 VDD P l=0.18u w=1.06u 
MM23 23 7 5 VDD P l=0.18u w=1.06u 
MM22 24 7 5 VDD P l=0.18u w=1.06u 
MM21 25 I1 VDD VDD P l=0.18u w=1.06u 
MM27 26 S1 28 VDD P l=0.18u w=1.06u 
MM20 26 S0 5 VDD P l=0.18u w=1.06u 
MM19 27 S0 5 VDD P l=0.18u w=1.06u 
MM18 VDD I0 28 VDD P l=0.187302u w=1.134u 
MM17 VDD S0 7 VDD P l=0.18u w=1.06u 
MM16 VDD S1 3 VDD P l=0.18u w=0.68u 
MM13 16 3 13 VSS N l=0.18u w=1u 
MM11 5 S0 13 VSS N l=0.18u w=1u 
MM12 14 S1 15 VSS N l=0.18u w=1u 
MM10 14 S0 5 VSS N l=0.18u w=1u 
MM9 Z 5 VSS VSS N l=0.18u w=0.58u 
MM8 15 I3 VSS VSS N l=0.18u w=1u 
MM7 VSS I1 16 VSS N l=0.18u w=1u 
MM6 5 7 17 VSS N l=0.185886u w=1.162u 
MM4 19 S1 17 VSS N l=0.18u w=1.01u 
MM5 5 7 18 VSS N l=0.18u w=1.1u 
MM14 18 3 20 VSS N l=0.18u w=1.1u 
MM15 VSS I2 19 VSS N l=0.186381u w=1.072u 
MM3 VSS I0 20 VSS N l=0.18u w=1.1u 
MM2 7 S0 VSS VSS N l=0.18u w=0.57u 
MM1 3 S1 VSS VSS N l=0.18u w=0.48u 
.ENDS mx04d0

.SUBCKT mx04d1 Z  I0 I1 I2 I3 S0 S1 VDD VSS
MM30 21 I2 VDD VDD P l=0.18u w=1.06u 
MM29 27 3 21 VDD P l=0.18u w=1.06u 
MM25 Z 5 VDD VDD P l=0.18u w=1.5u 
MM28 22 3 24 VDD P l=0.18u w=1.06u 
MM24 22 I3 VDD VDD P l=0.18u w=1.06u 
MM26 23 S1 25 VDD P l=0.18u w=1.06u 
MM23 23 7 5 VDD P l=0.18u w=1.06u 
MM22 24 7 5 VDD P l=0.18u w=1.06u 
MM21 25 I1 VDD VDD P l=0.18u w=1.06u 
MM27 26 S1 28 VDD P l=0.18u w=1.06u 
MM20 26 S0 5 VDD P l=0.18u w=1.06u 
MM19 27 S0 5 VDD P l=0.18u w=1.06u 
MM18 VDD I0 28 VDD P l=0.187302u w=1.134u 
MM17 VDD S0 7 VDD P l=0.18u w=1.06u 
MM16 VDD S1 3 VDD P l=0.18u w=0.68u 
MM13 16 3 13 VSS N l=0.18u w=1u 
MM11 5 S0 13 VSS N l=0.18u w=1u 
MM12 14 S1 15 VSS N l=0.18u w=1u 
MM10 14 S0 5 VSS N l=0.18u w=1u 
MM9 Z 5 VSS VSS N l=0.186381u w=1.072u 
MM8 15 I3 VSS VSS N l=0.18u w=1u 
MM7 VSS I1 16 VSS N l=0.18u w=1u 
MM6 5 7 17 VSS N l=0.185886u w=1.162u 
MM4 19 S1 17 VSS N l=0.18u w=1.01u 
MM5 5 7 18 VSS N l=0.18u w=1.1u 
MM14 18 3 20 VSS N l=0.18u w=1.1u 
MM15 VSS I2 19 VSS N l=0.186381u w=1.072u 
MM3 VSS I0 20 VSS N l=0.18u w=1.1u 
MM2 7 S0 VSS VSS N l=0.18u w=0.57u 
MM1 3 S1 VSS VSS N l=0.18u w=0.48u 
.ENDS mx04d1

.SUBCKT mx04d2 Z  I0 I1 I2 I3 S0 S1 VDD VSS
MM28 Z 4 VDD VDD P l=0.184379u w=1.562u 
MM27 Z 4 VDD VDD P l=0.18u w=1.5u 
MM31 21 2 23 VDD P l=0.18u w=1.06u 
MM26 21 I3 VDD VDD P l=0.18u w=1.06u 
MM29 22 S1 24 VDD P l=0.18u w=1.06u 
MM25 22 6 4 VDD P l=0.18u w=1.06u 
MM24 23 6 4 VDD P l=0.18u w=1.06u 
MM23 24 I1 VDD VDD P l=0.18u w=1.06u 
MM32 27 2 25 VDD P l=0.18u w=1.06u 
MM22 25 I2 VDD VDD P l=0.18u w=1.06u 
MM30 26 S1 28 VDD P l=0.18u w=1.06u 
MM21 26 S0 4 VDD P l=0.18u w=1.06u 
MM20 27 S0 4 VDD P l=0.18u w=1.06u 
MM19 VDD I0 28 VDD P l=0.187302u w=1.134u 
MM18 VDD S0 6 VDD P l=0.18u w=1.06u 
MM17 VDD S1 2 VDD P l=0.18u w=0.68u 
MM15 16 2 13 VSS N l=0.18u w=1.06u 
MM13 4 S0 13 VSS N l=0.18u w=1.06u 
MM14 14 S1 15 VSS N l=0.18u w=1.06u 
MM12 14 S0 4 VSS N l=0.18u w=1.06u 
MM11 Z 4 VSS VSS N l=0.187302u w=1.134u 
MM10 Z 4 VSS VSS N l=0.18u w=1.06u 
MM9 15 I3 VSS VSS N l=0.18u w=1.06u 
MM8 VSS I1 16 VSS N l=0.18u w=1.06u 
MM7 4 6 17 VSS N l=0.185886u w=1.162u 
MM5 19 S1 17 VSS N l=0.18u w=1.07u 
MM6 4 6 18 VSS N l=0.18u w=1.1u 
MM16 18 2 20 VSS N l=0.18u w=1.1u 
MM4 VSS I2 19 VSS N l=0.186042u w=1.132u 
MM3 VSS I0 20 VSS N l=0.18u w=1.1u 
MM2 6 S0 VSS VSS N l=0.18u w=0.57u 
MM1 2 S1 VSS VSS N l=0.18u w=0.48u 
.ENDS mx04d2

.SUBCKT mx04d4 Z  I0 I1 I2 I3 S0 S1 VDD VSS
MM35 23 S1 26 VDD P l=0.18u w=1.06u 
MM34 23 4 5 VDD P l=0.18u w=1.06u 
MM37 25 2 24 VDD P l=0.18u w=1.06u 
MM33 24 4 5 VDD P l=0.18u w=1.06u 
MM32 VDD 5 12 VDD P l=0.18u w=0.68u 
MM31 25 I3 VDD VDD P l=0.18u w=1.06u 
MM30 26 I1 VDD VDD P l=0.18u w=1.06u 
MM38 29 2 27 VDD P l=0.18u w=1.06u 
MM29 27 I2 VDD VDD P l=0.18u w=1.06u 
MM36 28 S1 30 VDD P l=0.18u w=1.06u 
MM28 28 S0 5 VDD P l=0.18u w=1.06u 
MM27 29 S0 5 VDD P l=0.18u w=1.06u 
MM26 VDD I0 30 VDD P l=0.187302u w=1.134u 
MM25 VDD S0 4 VDD P l=0.18u w=1.06u 
MM24 VDD 11 Z VDD P l=0.184906u w=1.59u 
MM23 VDD 11 Z VDD P l=0.18u w=1.52u 
MM22 Z 11 VDD VDD P l=0.18u w=1.52u 
MM21 VDD 12 11 VDD P l=0.184906u w=1.59u 
MM20 VDD S1 2 VDD P l=0.18u w=0.68u 
MM18 20 2 15 VSS N l=0.18u w=1u 
MM16 5 S0 15 VSS N l=0.18u w=1u 
MM17 16 S1 17 VSS N l=0.18u w=1u 
MM15 16 S0 5 VSS N l=0.18u w=1u 
MM14 12 5 VSS VSS N l=0.18u w=0.58u 
MM13 17 I3 VSS VSS N l=0.18u w=1u 
MM12 5 4 18 VSS N l=0.185886u w=1.162u 
MM10 21 S1 18 VSS N l=0.18u w=1.01u 
MM11 5 4 19 VSS N l=0.18u w=1.1u 
MM19 19 2 22 VSS N l=0.18u w=1.1u 
MM9 VSS I1 20 VSS N l=0.18u w=1u 
MM8 VSS I2 21 VSS N l=0.186381u w=1.072u 
MM7 VSS I0 22 VSS N l=0.18u w=1.1u 
MM6 4 S0 VSS VSS N l=0.18u w=0.57u 
MM4 Z 11 VSS VSS N l=0.186935u w=1.194u 
MM5 Z 11 VSS VSS N l=0.186935u w=1.194u 
MM3 Z 11 VSS VSS N l=0.18u w=1.12u 
MM2 VSS 12 11 VSS N l=0.18u w=1.12u 
MM1 2 S1 VSS VSS N l=0.18u w=0.48u 
.ENDS mx04d4

.SUBCKT nd02d0 ZN  A1 A2 VDD VSS
MM4 VDD A1 ZN VDD P l=0.18u w=0.94u 
MM3 VDD A2 ZN VDD P l=0.18u w=0.94u 
MM2 ZN A1 6 VSS N l=0.18u w=0.48u 
MM1 VSS A2 6 VSS N l=0.18u w=0.48u 
.ENDS nd02d0

.SUBCKT nd02d1 ZN  A1 A2 VDD VSS
MM4 ZN A1 VDD VDD P l=0.18u w=1.34u 
MM3 ZN A2 VDD VDD P l=0.18u w=1.34u 
MM2 ZN A1 6 VSS N l=0.18u w=0.82u 
MM1 VSS A2 6 VSS N l=0.18u w=0.82u 
.ENDS nd02d1

.SUBCKT nd02d2 ZN  A1 A2 VDD VSS
MM7 ZN A1 VDD VDD P l=0.18u w=1.32u 
MM6 VDD A2 ZN VDD P l=0.186913u w=1.406u 
MM8 ZN A1 VDD VDD P l=0.186591u w=1.402u 
MM5 VDD A2 ZN VDD P l=0.18u w=1.32u 
MM4 7 A1 ZN VSS N l=0.18u w=0.9u 
MM3 6 A1 ZN VSS N l=0.18u w=0.9u 
MM2 6 A2 VSS VSS N l=0.18u w=0.9u 
MM1 7 A2 VSS VSS N l=0.18u w=0.9u 
.ENDS nd02d2

.SUBCKT nd02d4 ZN  A1 A2 VDD VSS
MM12 VDD 2 3 VDD P l=0.185597u w=1.222u 
MM10 ZN 3 VDD VDD P l=0.183417u w=2.002u 
MM11 VDD 3 ZN VDD P l=0.183417u w=2.002u 
MM9 VDD 3 ZN VDD P l=0.183417u w=2.002u 
MM8 VDD A1 2 VDD P l=0.18u w=0.94u 
MM7 VDD A2 2 VDD P l=0.186826u w=1.002u 
MM6 3 2 VSS VSS N l=0.186381u w=1.072u 
MM5 ZN 3 VSS VSS N l=0.185135u w=1.332u 
MM4 ZN 3 VSS VSS N l=0.185135u w=1.332u 
MM3 ZN 3 VSS VSS N l=0.185135u w=1.332u 
MM2 8 A1 2 VSS N l=0.18u w=0.48u 
MM1 8 A2 VSS VSS N l=0.18u w=0.48u 
.ENDS nd02d4

.SUBCKT nd03d0 ZN  A1 A2 A3 VDD VSS
MM6 VDD A2 ZN VDD P l=0.18u w=0.52u 
MM5 ZN A1 VDD VDD P l=0.18u w=0.52u 
MM4 VDD A3 ZN VDD P l=0.18u w=0.52u 
MM3 7 A2 8 VSS N l=0.18u w=0.48u 
MM2 VSS A1 7 VSS N l=0.18u w=0.48u 
MM1 ZN A3 8 VSS N l=0.18u w=0.48u 
.ENDS nd03d0

.SUBCKT nd03d1 ZN  A1 A2 A3 VDD VSS
MM6 VDD A2 ZN VDD P l=0.185059u w=1.352u 
MM5 VDD A1 ZN VDD P l=0.18607u w=1.364u 
MM4 VDD A3 ZN VDD P l=0.185692u w=1.286u 
MM2 7 A1 ZN VSS N l=0.18u w=1.09u 
MM3 8 A2 7 VSS N l=0.18u w=1.09u 
MM1 8 A3 VSS VSS N l=0.185937u w=1.152u 
.ENDS nd03d1

.SUBCKT nd03d2 ZN  A1 A2 A3 VDD VSS
MM12 VDD A3 ZN VDD P l=0.185006u w=1.654u 
MM11 VDD A3 ZN VDD P l=0.18u w=1.58u 
MM10 VDD A1 ZN VDD P l=0.191693u w=1.565u 
MM9 VDD A1 ZN VDD P l=0.184166u w=1.642u 
MM8 ZN A2 VDD VDD P l=0.184727u w=1.65u 
MM7 ZN A2 VDD VDD P l=0.18u w=1.58u 
MM6 ZN A3 9 VSS N l=0.18u w=1.09u 
MM5 ZN A3 8 VSS N l=0.18u w=1.09u 
MM4 VSS A1 7 VSS N l=0.186264u w=1.092u 
MM2 8 A2 7 VSS N l=0.18u w=1.09u 
MM1 9 A2 10 VSS N l=0.18u w=1.09u 
MM3 VSS A1 10 VSS N l=0.18u w=1.09u 
.ENDS nd03d2

.SUBCKT nd03d4 ZN  A1 A2 A3 VDD VSS
MM14 3 2 VDD VDD P l=0.185253u w=1.302u 
MM12 VDD 3 ZN VDD P l=0.183417u w=2.002u 
MM13 VDD 3 ZN VDD P l=0.183417u w=2.002u 
MM11 VDD 3 ZN VDD P l=0.183417u w=2.002u 
MM10 2 A3 VDD VDD P l=0.18u w=0.52u 
MM9 2 A2 VDD VDD P l=0.18u w=0.52u 
MM8 2 A1 VDD VDD P l=0.18u w=0.52u 
MM7 VSS 2 3 VSS N l=0.186381u w=1.072u 
MM6 ZN 3 VSS VSS N l=0.185135u w=1.332u 
MM5 ZN 3 VSS VSS N l=0.185135u w=1.332u 
MM4 VSS 3 ZN VSS N l=0.185135u w=1.332u 
MM3 2 A3 9 VSS N l=0.18u w=0.48u 
MM2 10 A2 9 VSS N l=0.18u w=0.48u 
MM1 VSS A1 10 VSS N l=0.18u w=0.48u 
.ENDS nd03d4

.SUBCKT nd04d0 ZN  A1 A2 A3 A4 VDD VSS
MM8 VDD A2 ZN VDD P l=0.18u w=0.63u 
MM7 VDD A3 ZN VDD P l=0.18u w=0.63u 
MM6 VDD A1 ZN VDD P l=0.18u w=0.63u 
MM5 VDD A4 ZN VDD P l=0.18u w=0.63u 
MM4 8 A2 ZN VSS N l=0.18u w=0.6u 
MM3 8 A3 9 VSS N l=0.18u w=0.6u 
MM2 10 A1 9 VSS N l=0.18u w=0.6u 
MM1 10 A4 VSS VSS N l=0.18u w=0.6u 
.ENDS nd04d0

.SUBCKT nd04d1 ZN  A1 A2 A3 A4 VDD VSS
MM8 VDD A3 ZN VDD P l=0.185691u w=1.202u 
MM7 ZN A2 VDD VDD P l=0.18u w=1.2u 
MM6 ZN A1 VDD VDD P l=0.185691u w=1.202u 
MM5 VDD A4 ZN VDD P l=0.18u w=1.2u 
MM3 ZN A2 8 VSS N l=0.18u w=1.11u 
MM4 8 A3 9 VSS N l=0.18u w=1.11u 
MM2 10 A1 9 VSS N l=0.18u w=1.11u 
MM1 10 A4 VSS VSS N l=0.18u w=1.11u 
.ENDS nd04d1

.SUBCKT nd04d2 ZN  A1 A2 A3 A4 VDD VSS
MM14 VDD A3 6 VDD P l=0.185691u w=1.202u 
MM12 VDD A2 6 VDD P l=0.18u w=1.2u 
MM13 6 A1 VDD VDD P l=0.185691u w=1.202u 
MM11 VDD A4 6 VDD P l=0.18u w=1.2u 
MM10 7 6 VDD VDD P l=0.185253u w=1.302u 
MM9 VDD 7 ZN VDD P l=0.184554u w=1.502u 
MM8 ZN 7 VDD VDD P l=0.184554u w=1.502u 
MM5 6 A2 11 VSS N l=0.18u w=1.11u 
MM7 10 A3 11 VSS N l=0.18u w=1.11u 
MM6 12 A1 10 VSS N l=0.18u w=1.11u 
MM4 12 A4 VSS VSS N l=0.18u w=1.11u 
MM3 VSS 6 7 VSS N l=0.186381u w=1.072u 
MM2 VSS 7 ZN VSS N l=0.186826u w=1.002u 
MM1 VSS 7 ZN VSS N l=0.186826u w=1.002u 
.ENDS nd04d2

.SUBCKT nd04d4 ZN  A1 A2 A3 A4 VDD VSS
MM16 VDD A3 6 VDD P l=0.185691u w=1.202u 
MM14 VDD A2 6 VDD P l=0.18u w=1.2u 
MM15 6 A1 VDD VDD P l=0.185691u w=1.202u 
MM13 VDD A4 6 VDD P l=0.18u w=1.2u 
MM12 7 6 VDD VDD P l=0.185253u w=1.302u 
MM10 VDD 7 ZN VDD P l=0.183417u w=2.002u 
MM11 ZN 7 VDD VDD P l=0.183417u w=2.002u 
MM9 ZN 7 VDD VDD P l=0.183417u w=2.002u 
MM8 VSS 6 7 VSS N l=0.186381u w=1.072u 
MM7 ZN 7 VSS VSS N l=0.185135u w=1.332u 
MM6 VSS 7 ZN VSS N l=0.185135u w=1.332u 
MM5 VSS 7 ZN VSS N l=0.185135u w=1.332u 
MM2 6 A2 11 VSS N l=0.18u w=1.11u 
MM4 10 A3 11 VSS N l=0.18u w=1.11u 
MM3 12 A1 10 VSS N l=0.18u w=1.11u 
MM1 12 A4 VSS VSS N l=0.18u w=1.11u 
.ENDS nd04d4

.SUBCKT nd12d0 ZN  A1 A2 VDD VSS
MM6 VDD 2 ZN VDD P l=0.18u w=0.62u 
MM5 VDD A2 ZN VDD P l=0.18u w=0.62u 
MM4 VDD A1 2 VDD P l=0.18u w=0.62u 
MM2 ZN A2 7 VSS N l=0.18u w=0.48u 
MM3 VSS 2 7 VSS N l=0.18u w=0.48u 
MM1 VSS A1 2 VSS N l=0.18u w=0.48u 
.ENDS nd12d0

.SUBCKT nd12d1 ZN  A1 A2 VDD VSS
MM6 VDD 2 ZN VDD P l=0.184554u w=1.502u 
MM5 VDD A2 ZN VDD P l=0.184554u w=1.502u 
MM4 VDD A1 2 VDD P l=0.186618u w=1.106u 
MM3 7 2 VSS VSS N l=0.189184u w=1.091u 
MM2 7 A2 ZN VSS N l=0.18u w=1u 
MM1 VSS A1 2 VSS N l=0.18u w=0.57u 
.ENDS nd12d1

.SUBCKT nd12d2 ZN  A1 A2 VDD VSS
MM9 ZN A2 VDD VDD P l=0.18u w=1.54u 
MM8 ZN 3 VDD VDD P l=0.18513u w=1.614u 
MM10 VDD A2 ZN VDD P l=0.18u w=1.54u 
MM7 VDD 3 ZN VDD P l=0.18u w=1.54u 
MM6 VDD A1 3 VDD P l=0.184558u w=1.606u 
MM5 ZN A2 7 VSS N l=0.18u w=1.03u 
MM4 ZN A2 8 VSS N l=0.18u w=1.03u 
MM3 VSS 3 7 VSS N l=0.190885u w=1.141u 
MM2 VSS 3 8 VSS N l=0.18u w=1.03u 
MM1 3 A1 VSS VSS N l=0.18u w=1.03u 
.ENDS nd12d2

.SUBCKT nd12d4 ZN  A1 A2 VDD VSS
MM14 3 2 VDD VDD P l=0.185597u w=1.222u 
MM12 VDD 3 ZN VDD P l=0.183417u w=2.002u 
MM13 VDD 3 ZN VDD P l=0.183417u w=2.002u 
MM11 ZN 3 VDD VDD P l=0.183417u w=2.002u 
MM10 VDD A1 6 VDD P l=0.18u w=1.11u 
MM9 VDD A2 2 VDD P l=0.184615u w=1.482u 
MM8 VDD 6 2 VDD P l=0.184615u w=1.482u 
MM7 VSS 2 3 VSS N l=0.186381u w=1.072u 
MM6 VSS 3 ZN VSS N l=0.185135u w=1.332u 
MM5 VSS 3 ZN VSS N l=0.185135u w=1.332u 
MM4 VSS 3 ZN VSS N l=0.185135u w=1.332u 
MM3 VSS A1 6 VSS N l=0.18u w=0.57u 
MM2 2 A2 9 VSS N l=0.18u w=1u 
MM1 9 6 VSS VSS N l=0.189184u w=1.091u 
.ENDS nd12d4

.SUBCKT nd13d1 ZN  A1 A2 A3 VDD VSS
MM7 ZN A2 VDD VDD P l=0.184949u w=1.382u 
MM8 VDD A3 ZN VDD P l=0.184949u w=1.382u 
MM6 VDD 4 ZN VDD P l=0.184949u w=1.382u 
MM5 VDD A1 4 VDD P l=0.185281u w=1.386u 
MM3 8 A2 ZN VSS N l=0.18u w=1.01u 
MM4 9 A3 8 VSS N l=0.18u w=1.01u 
MM2 9 4 VSS VSS N l=0.18u w=1.01u 
MM1 4 A1 VSS VSS N l=0.187091u w=1.1u 
.ENDS nd13d1

.SUBCKT nd13d2 ZN  A1 A2 A3 VDD VSS
MM14 VDD A3 ZN VDD P l=0.185067u w=1.634u 
MM13 ZN A3 VDD VDD P l=0.18u w=1.56u 
MM12 VDD A2 ZN VDD P l=0.184217u w=1.622u 
MM11 VDD A2 ZN VDD P l=0.18u w=1.56u 
MM10 ZN 4 VDD VDD P l=0.184217u w=1.622u 
MM9 ZN 4 VDD VDD P l=0.18u w=1.56u 
MM8 VDD A1 4 VDD P l=0.18u w=0.7u 
MM7 9 A3 ZN VSS N l=0.186207u w=1.102u 
MM6 8 A3 ZN VSS N l=0.186207u w=1.102u 
MM5 11 A2 8 VSS N l=0.18u w=1.04u 
MM4 10 A2 9 VSS N l=0.18u w=1.04u 
MM3 10 4 VSS VSS N l=0.18u w=1.04u 
MM2 11 4 VSS VSS N l=0.18u w=1.04u 
MM1 VSS A1 4 VSS N l=0.18u w=0.72u 
.ENDS nd13d2

.SUBCKT nd13d4 ZN  A1 A2 A3 VDD VSS
MM16 6 A2 VDD VDD P l=0.184949u w=1.382u 
MM15 VDD A3 6 VDD P l=0.184949u w=1.382u 
MM14 VDD 4 6 VDD P l=0.184949u w=1.382u 
MM13 VDD A1 4 VDD P l=0.185281u w=1.386u 
MM12 7 6 VDD VDD P l=0.185597u w=1.222u 
MM10 ZN 7 VDD VDD P l=0.183417u w=2.002u 
MM11 ZN 7 VDD VDD P l=0.183417u w=2.002u 
MM9 ZN 7 VDD VDD P l=0.183417u w=2.002u 
MM8 7 6 VSS VSS N l=0.186381u w=1.072u 
MM7 ZN 7 VSS VSS N l=0.185135u w=1.332u 
MM6 ZN 7 VSS VSS N l=0.185135u w=1.332u 
MM5 ZN 7 VSS VSS N l=0.185135u w=1.332u 
MM4 10 A2 6 VSS N l=0.18u w=1.01u 
MM3 11 A3 10 VSS N l=0.18u w=1.01u 
MM2 11 4 VSS VSS N l=0.18u w=1.01u 
MM1 4 A1 VSS VSS N l=0.187091u w=1.1u 
.ENDS nd13d4

.SUBCKT nd23d1 ZN  A1 A2 A3 VDD VSS
MM10 VDD A2 6 VDD P l=0.18u w=0.59u 
MM9 VDD A1 4 VDD P l=0.18u w=0.59u 
MM8 VDD 4 ZN VDD P l=0.184674u w=1.566u 
MM7 ZN A3 VDD VDD P l=0.184968u w=1.57u 
MM6 VDD 6 ZN VDD P l=0.18u w=1.5u 
MM5 ZN 4 10 VSS N l=0.18u w=1.11u 
MM4 VSS A3 9 VSS N l=0.18u w=1.11u 
MM3 9 6 10 VSS N l=0.18u w=1.11u 
MM2 6 A2 VSS VSS N l=0.18u w=0.66u 
MM1 VSS A1 4 VSS N l=0.18u w=0.48u 
.ENDS nd23d1

.SUBCKT nd23d2 ZN  A1 A2 A3 VDD VSS
MM12 VDD 2 ZN VDD P l=0.18u w=1.5u 
MM11 VDD 2 ZN VDD P l=0.18u w=1.5u 
MM10 9 A1 VDD VDD P l=0.18u w=1.19u 
MM9 9 A2 10 VDD P l=0.18u w=1.19u 
MM8 2 5 10 VDD P l=0.18u w=1.19u 
MM7 VDD A3 5 VDD P l=0.18u w=0.51u 
MM6 ZN 2 VSS VSS N l=0.18u w=1u 
MM5 ZN 2 VSS VSS N l=0.18u w=1u 
MM4 VSS A1 2 VSS N l=0.18u w=0.48u 
MM3 VSS A2 2 VSS N l=0.18u w=0.48u 
MM2 VSS 5 2 VSS N l=0.18u w=0.48u 
MM1 VSS A3 5 VSS N l=0.18u w=0.49u 
.ENDS nd23d2

.SUBCKT nd23d4 ZN  A1 A2 A3 VDD VSS
MM13 ZN 3 VDD VDD P l=0.183881u w=2.01u 
MM12 VDD 3 ZN VDD P l=0.18516u w=2.035u 
MM11 VDD 3 ZN VDD P l=0.18u w=1.94u 
MM14 9 A1 VDD VDD P l=0.18u w=1.19u 
MM10 9 A2 10 VDD P l=0.18u w=1.19u 
MM9 3 5 10 VDD P l=0.18u w=1.19u 
MM8 VDD A3 5 VDD P l=0.18u w=0.51u 
MM6 ZN 3 VSS VSS N l=0.187962u w=1.379u 
MM5 ZN 3 VSS VSS N l=0.185097u w=1.342u 
MM4 ZN 3 VSS VSS N l=0.18u w=1.28u 
MM7 VSS A1 3 VSS N l=0.18u w=0.48u 
MM3 VSS A2 3 VSS N l=0.18u w=0.48u 
MM2 VSS 5 3 VSS N l=0.18u w=0.48u 
MM1 VSS A3 5 VSS N l=0.18u w=0.49u 
.ENDS nd23d4

.SUBCKT nr02d0 ZN  A1 A2 VDD VSS
MM4 VDD A2 6 VDD P l=0.18u w=0.89u 
MM3 ZN A1 6 VDD P l=0.18u w=0.89u 
MM2 VSS A2 ZN VSS N l=0.18u w=0.48u 
MM1 ZN A1 VSS VSS N l=0.18u w=0.48u 
.ENDS nr02d0

.SUBCKT nr02d1 ZN  A1 A2 VDD VSS
MM3 6 A2 ZN VDD P l=0.186659u w=1.649u 
MM4 6 A1 VDD VDD P l=0.186659u w=1.649u 
MM2 VSS A1 ZN VSS N l=0.18u w=0.89u 
MM1 VSS A2 ZN VSS N l=0.18u w=0.89u 
.ENDS nr02d1

.SUBCKT nr02d2 ZN  A1 A2 VDD VSS
MM8 6 A1 ZN VDD P l=0.187294u w=1.637u 
MM7 ZN A1 7 VDD P l=0.18u w=1.53u 
MM6 6 A2 VDD VDD P l=0.188u w=1.65u 
MM5 VDD A2 7 VDD P l=0.186015u w=1.616u 
MM4 VSS A1 ZN VSS N l=0.188861u w=1.185u 
MM3 VSS A1 ZN VSS N l=0.18u w=1.09u 
MM2 ZN A2 VSS VSS N l=0.186724u w=1.16u 
MM1 ZN A2 VSS VSS N l=0.18u w=1.09u 
.ENDS nr02d2

.SUBCKT nr02d4 ZN  A1 A2 VDD VSS
MM12 VDD 2 3 VDD P l=0.185022u w=1.362u 
MM11 VDD 3 ZN VDD P l=0.184682u w=2.076u 
MM10 VDD 3 ZN VDD P l=0.18u w=1.99u 
MM9 ZN 3 VDD VDD P l=0.18u w=1.99u 
MM8 VDD A1 8 VDD P l=0.18u w=0.75u 
MM7 8 A2 2 VDD P l=0.18u w=0.75u 
MM6 3 2 VSS VSS N l=0.18u w=0.86u 
MM4 ZN 3 VSS VSS N l=0.185294u w=1.564u 
MM5 ZN 3 VSS VSS N l=0.186168u w=1.576u 
MM3 ZN 3 VSS VSS N l=0.18u w=1.49u 
MM2 VSS A1 2 VSS N l=0.18u w=0.5u 
MM1 VSS A2 2 VSS N l=0.18u w=0.5u 
.ENDS nr02d4

.SUBCKT nr03d0 ZN  A1 A2 A3 VDD VSS
MM6 8 A2 7 VDD P l=0.18u w=0.8u 
MM5 VDD A1 7 VDD P l=0.18u w=0.8u 
MM4 8 A3 ZN VDD P l=0.18u w=0.8u 
MM3 VSS A2 ZN VSS N l=0.18u w=0.52u 
MM2 VSS A1 ZN VSS N l=0.18u w=0.52u 
MM1 ZN A3 VSS VSS N l=0.18u w=0.52u 
.ENDS nr03d0

.SUBCKT nr03d1 ZN  A1 A2 A3 VDD VSS
MM6 8 A2 7 VDD P l=0.18u w=1.32u 
MM5 7 A1 VDD VDD P l=0.188679u w=1.431u 
MM4 8 A3 ZN VDD P l=0.18u w=1.32u 
MM3 VSS A2 ZN VSS N l=0.18u w=1.14u 
MM2 VSS A1 ZN VSS N l=0.18u w=0.85u 
MM1 VSS A3 ZN VSS N l=0.18814u w=1.231u 
.ENDS nr03d1

.SUBCKT nr03d2 ZN  A1 A2 A3 VDD VSS
MM12 3 2 VDD VDD P l=0.185097u w=1.342u 
MM11 ZN 3 VDD VDD P l=0.184554u w=1.502u 
MM10 VDD 3 ZN VDD P l=0.184861u w=1.506u 
MM9 9 A3 VDD VDD P l=0.185925u w=1.691u 
MM8 10 A2 9 VDD P l=0.18u w=1.6u 
MM7 10 A1 2 VDD P l=0.18u w=1.6u 
MM6 VSS 2 3 VSS N l=0.186381u w=1.072u 
MM5 ZN 3 VSS VSS N l=0.187276u w=1.006u 
MM4 VSS 3 ZN VSS N l=0.186826u w=1.002u 
MM3 VSS A3 2 VSS N l=0.185989u w=1.142u 
MM2 VSS A2 2 VSS N l=0.18u w=1.08u 
MM1 2 A1 VSS VSS N l=0.186387u w=1.146u 
.ENDS nr03d2

.SUBCKT nr03d4 ZN  A1 A2 A3 VDD VSS
MM14 3 2 VDD VDD P l=0.184985u w=1.372u 
MM13 VDD 3 ZN VDD P l=0.183881u w=2.01u 
MM12 VDD 3 ZN VDD P l=0.18516u w=2.035u 
MM11 ZN 3 VDD VDD P l=0.18u w=1.94u 
MM10 9 A3 VDD VDD P l=0.185925u w=1.691u 
MM9 10 A2 9 VDD P l=0.18u w=1.6u 
MM8 10 A1 2 VDD P l=0.18u w=1.6u 
MM7 VSS 2 3 VSS N l=0.186867u w=1.066u 
MM6 ZN 3 VSS VSS N l=0.188286u w=1.383u 
MM5 VSS 3 ZN VSS N l=0.185097u w=1.342u 
MM4 ZN 3 VSS VSS N l=0.18u w=1.28u 
MM3 VSS A3 2 VSS N l=0.185989u w=1.142u 
MM2 VSS A2 2 VSS N l=0.18u w=1.08u 
MM1 2 A1 VSS VSS N l=0.186387u w=1.146u 
.ENDS nr03d4

.SUBCKT nr04d0 ZN  A1 A2 A3 A4 VDD VSS
MM8 VDD A1 8 VDD P l=0.18u w=0.87u 
MM7 9 A2 8 VDD P l=0.18u w=0.87u 
MM6 9 A3 10 VDD P l=0.18u w=0.87u 
MM5 ZN A4 10 VDD P l=0.18u w=0.87u 
MM4 ZN A1 VSS VSS N l=0.18u w=0.48u 
MM3 VSS A2 ZN VSS N l=0.18u w=0.48u 
MM2 ZN A3 VSS VSS N l=0.18u w=0.48u 
MM1 ZN A4 VSS VSS N l=0.18u w=0.48u 
.ENDS nr04d0

.SUBCKT nr04d1 ZN  A1 A2 A3 A4 VDD VSS
MM7 9 A2 8 VDD P l=0.18u w=1.55u 
MM6 8 A3 10 VDD P l=0.18481u w=1.422u 
MM8 9 A1 VDD VDD P l=0.18u w=1.55u 
MM5 ZN A4 10 VDD P l=0.18481u w=1.422u 
MM4 VSS A1 ZN VSS N l=0.18u w=0.96u 
MM3 ZN A2 VSS VSS N l=0.18u w=0.96u 
MM2 ZN A3 VSS VSS N l=0.18u w=0.89u 
MM1 ZN A4 VSS VSS N l=0.18u w=0.89u 
.ENDS nr04d1

.SUBCKT nr04d2 ZN  A1 A2 A3 A4 VDD VSS
MM13 6 A1 10 VDD P l=0.18481u w=1.422u 
MM14 11 A2 10 VDD P l=0.18481u w=1.422u 
MM11 12 A3 11 VDD P l=0.18u w=1.55u 
MM12 12 A4 VDD VDD P l=0.18u w=1.55u 
MM10 7 6 VDD VDD P l=0.185097u w=1.342u 
MM9 ZN 7 VDD VDD P l=0.184554u w=1.502u 
MM8 VDD 7 ZN VDD P l=0.184861u w=1.506u 
MM7 6 A2 VSS VSS N l=0.18u w=0.89u 
MM6 6 A1 VSS VSS N l=0.18u w=0.89u 
MM5 VSS A4 6 VSS N l=0.18u w=0.96u 
MM4 6 A3 VSS VSS N l=0.18u w=0.96u 
MM3 VSS 6 7 VSS N l=0.186381u w=1.072u 
MM2 ZN 7 VSS VSS N l=0.187276u w=1.006u 
MM1 VSS 7 ZN VSS N l=0.186826u w=1.002u 
.ENDS nr04d2

.SUBCKT nr04d4 ZN  A1 A2 A3 A4 VDD VSS
MM16 3 2 VDD VDD P l=0.18532u w=1.376u 
MM15 VDD 3 ZN VDD P l=0.183881u w=2.01u 
MM14 ZN 3 VDD VDD P l=0.18516u w=2.035u 
MM13 ZN 3 VDD VDD P l=0.18u w=1.94u 
MM11 2 A1 10 VDD P l=0.18481u w=1.422u 
MM12 11 A2 10 VDD P l=0.18481u w=1.422u 
MM9 12 A3 11 VDD P l=0.18u w=1.55u 
MM10 12 A4 VDD VDD P l=0.18u w=1.55u 
MM8 VSS 2 3 VSS N l=0.186441u w=1.062u 
MM7 ZN 3 VSS VSS N l=0.187636u w=1.375u 
MM6 VSS 3 ZN VSS N l=0.185438u w=1.346u 
MM5 VSS 3 ZN VSS N l=0.18u w=1.28u 
MM4 VSS A2 2 VSS N l=0.18u w=0.89u 
MM3 2 A1 VSS VSS N l=0.18u w=0.89u 
MM2 VSS A4 2 VSS N l=0.18u w=0.96u 
MM1 2 A3 VSS VSS N l=0.18u w=0.96u 
.ENDS nr04d4

.SUBCKT nr13d1 ZN  A1 A2 A3 VDD VSS
MM8 ZN A3 8 VDD P l=0.18u w=1.91u 
MM7 8 A2 9 VDD P l=0.18u w=1.91u 
MM6 VDD A1 5 VDD P l=0.18u w=0.82u 
MM5 VDD 5 9 VDD P l=0.18u w=1.91u 
MM4 ZN A3 VSS VSS N l=0.18532u w=1.376u 
MM2 VSS A1 5 VSS N l=0.18u w=0.5u 
MM3 ZN A2 VSS VSS N l=0.184985u w=1.372u 
MM1 ZN 5 VSS VSS N l=0.184985u w=1.372u 
.ENDS nr13d1

.SUBCKT nr13d2 ZN  A1 A2 A3 VDD VSS
MM14 VDD 2 7 VDD P l=0.186094u w=1.28u 
MM13 5 A2 VDD VDD P l=0.18u w=0.97u 
MM12 VDD A1 7 VDD P l=0.185737u w=1.276u 
MM11 VDD 5 7 VDD P l=0.188388u w=1.309u 
MM10 VDD A3 2 VDD P l=0.18u w=0.5u 
MM9 VDD 7 ZN VDD P l=0.185398u w=1.534u 
MM8 VDD 7 ZN VDD P l=0.18u w=1.46u 
MM7 VSS A3 2 VSS N l=0.18u w=0.48u 
MM6 VSS 7 ZN VSS N l=0.18u w=1u 
MM5 VSS 7 ZN VSS N l=0.18u w=1u 
MM4 7 2 10 VSS N l=0.18u w=1.49u 
MM3 VSS A2 5 VSS N l=0.18u w=0.61u 
MM2 11 A1 10 VSS N l=0.18u w=1.49u 
MM1 VSS 5 11 VSS N l=0.18u w=1.49u 
.ENDS nr13d2

.SUBCKT nr13d4 ZN  A1 A2 A3 VDD VSS
MM16 4 A2 VDD VDD P l=0.18u w=0.97u 
MM15 VDD A1 7 VDD P l=0.185377u w=1.272u 
MM14 VDD 4 7 VDD P l=0.185213u w=1.312u 
MM13 7 5 VDD VDD P l=0.18u w=1.28u 
MM12 VDD A3 5 VDD P l=0.18u w=0.5u 
MM10 VDD 7 ZN VDD P l=0.184091u w=2.024u 
MM11 ZN 7 VDD VDD P l=0.184091u w=2.024u 
MM9 ZN 7 VDD VDD P l=0.18u w=1.95u 
MM8 VSS A3 5 VSS N l=0.18u w=0.59u 
MM7 VSS 7 ZN VSS N l=0.18u w=1.33u 
MM6 VSS 7 ZN VSS N l=0.18u w=1.33u 
MM5 ZN 7 VSS VSS N l=0.18u w=1.33u 
MM4 VSS A2 4 VSS N l=0.18u w=0.61u 
MM3 10 A1 11 VSS N l=0.18u w=1.49u 
MM2 VSS 4 10 VSS N l=0.18u w=1.49u 
MM1 7 5 11 VSS N l=0.18u w=1.49u 
.ENDS nr13d4

.SUBCKT nr23d1 ZN  A1 A2 A3 VDD VSS
MM10 3 A2 VDD VDD P l=0.18u w=0.5u 
MM9 ZN 3 9 VDD P l=0.18u w=1.88u 
MM8 VDD A1 6 VDD P l=0.18u w=0.5u 
MM7 10 A3 9 VDD P l=0.18u w=1.88u 
MM6 VDD 6 10 VDD P l=0.18u w=1.88u 
MM5 VSS 3 ZN VSS N l=0.189333u w=1.125u 
MM4 VSS A1 6 VSS N l=0.18u w=0.48u 
MM3 VSS A3 ZN VSS N l=0.18u w=1.02u 
MM2 ZN 6 VSS VSS N l=0.187156u w=1.09u 
MM1 3 A2 VSS VSS N l=0.18u w=0.49u 
.ENDS nr23d1

.SUBCKT nr23d2 ZN  A1 A2 A3 VDD VSS
MM12 VDD A3 4 VDD P l=0.18u w=0.54u 
MM11 ZN 3 VDD VDD P l=0.18u w=1.5u 
MM10 VDD 3 ZN VDD P l=0.18u w=1.5u 
MM9 3 4 VDD VDD P l=0.185692u w=1.286u 
MM8 3 A2 VDD VDD P l=0.185335u w=1.282u 
MM7 VDD A1 3 VDD P l=0.186047u w=1.29u 
MM6 VSS A3 4 VSS N l=0.18u w=0.48u 
MM5 ZN 3 VSS VSS N l=0.18u w=1u 
MM4 ZN 3 VSS VSS N l=0.18u w=1u 
MM3 9 4 3 VSS N l=0.18u w=1.49u 
MM2 10 A2 9 VSS N l=0.18u w=1.49u 
MM1 10 A1 VSS VSS N l=0.18u w=1.49u 
.ENDS nr23d2

.SUBCKT nr23d4 ZN  A1 A2 A3 VDD VSS
MM14 VDD A3 4 VDD P l=0.18u w=0.54u 
MM13 VDD 3 ZN VDD P l=0.183881u w=2.01u 
MM12 VDD 3 ZN VDD P l=0.18516u w=2.035u 
MM11 VDD 3 ZN VDD P l=0.18u w=1.94u 
MM10 3 4 VDD VDD P l=0.185692u w=1.286u 
MM9 3 A2 VDD VDD P l=0.185335u w=1.282u 
MM8 VDD A1 3 VDD P l=0.186047u w=1.29u 
MM7 VSS A3 4 VSS N l=0.18u w=0.48u 
MM6 ZN 3 VSS VSS N l=0.188286u w=1.383u 
MM5 VSS 3 ZN VSS N l=0.185097u w=1.342u 
MM4 ZN 3 VSS VSS N l=0.18u w=1.28u 
MM3 9 4 3 VSS N l=0.18u w=1.49u 
MM2 10 A2 9 VSS N l=0.18u w=1.49u 
MM1 10 A1 VSS VSS N l=0.18u w=1.49u 
.ENDS nr23d4

.SUBCKT oai211d1 ZN  A B C1 C2 VDD VSS
MM8 ZN A VDD VDD P l=0.185692u w=1.286u 
MM7 ZN B VDD VDD P l=0.18u w=1.37u 
MM6 10 C1 ZN VDD P l=0.183333u w=2.052u 
MM5 10 C2 VDD VDD P l=0.18356u w=2.056u 
MM4 ZN A 9 VSS N l=0.18u w=1.14u 
MM3 9 B 8 VSS N l=0.18u w=1.14u 
MM2 VSS C1 8 VSS N l=0.185691u w=1.202u 
MM1 8 C2 VSS VSS N l=0.187156u w=1.09u 
.ENDS oai211d1

.SUBCKT oai211d2 ZN  A B C1 C2 VDD VSS
MM14 6 A VDD VDD P l=0.18u w=1.31u 
MM13 6 B VDD VDD P l=0.184985u w=1.372u 
MM12 12 C1 6 VDD P l=0.183333u w=2.052u 
MM11 12 C2 VDD VDD P l=0.18356u w=2.056u 
MM10 7 6 VDD VDD P l=0.185597u w=1.222u 
MM9 VDD 7 ZN VDD P l=0.184554u w=1.502u 
MM8 ZN 7 VDD VDD P l=0.184554u w=1.502u 
MM7 6 A 11 VSS N l=0.18u w=1.14u 
MM6 11 B 10 VSS N l=0.18u w=1.14u 
MM5 VSS C1 10 VSS N l=0.185691u w=1.202u 
MM4 10 C2 VSS VSS N l=0.187156u w=1.09u 
MM3 VSS 6 7 VSS N l=0.186381u w=1.072u 
MM2 VSS 7 ZN VSS N l=0.186826u w=1.002u 
MM1 VSS 7 ZN VSS N l=0.186826u w=1.002u 
.ENDS oai211d2

.SUBCKT oai211d4 ZN  A B C1 C2 VDD VSS
MM16 3 2 VDD VDD P l=0.185597u w=1.222u 
MM14 VDD 3 ZN VDD P l=0.183417u w=2.002u 
MM15 ZN 3 VDD VDD P l=0.183417u w=2.002u 
MM13 ZN 3 VDD VDD P l=0.183417u w=2.002u 
MM12 2 A VDD VDD P l=0.185562u w=1.316u 
MM11 2 B VDD VDD P l=0.18u w=1.37u 
MM10 12 C1 2 VDD P l=0.183333u w=2.052u 
MM9 12 C2 VDD VDD P l=0.18356u w=2.056u 
MM8 VSS 2 3 VSS N l=0.186381u w=1.072u 
MM7 ZN 3 VSS VSS N l=0.185135u w=1.332u 
MM6 VSS 3 ZN VSS N l=0.185135u w=1.332u 
MM5 VSS 3 ZN VSS N l=0.185135u w=1.332u 
MM4 2 A 11 VSS N l=0.18u w=1.14u 
MM3 11 B 10 VSS N l=0.18u w=1.14u 
MM2 VSS C1 10 VSS N l=0.185691u w=1.202u 
MM1 10 C2 VSS VSS N l=0.187156u w=1.09u 
.ENDS oai211d4

.SUBCKT oai21d1 ZN  A B1 B2 VDD VSS
MM6 8 B1 ZN VDD P l=0.18u w=1.31u 
MM5 VDD A ZN VDD P l=0.185213u w=1.312u 
MM4 8 B2 VDD VDD P l=0.18u w=1.31u 
MM3 VSS B1 6 VSS N l=0.186441u w=1.062u 
MM2 ZN A 6 VSS N l=0.18u w=1.09u 
MM1 6 B2 VSS VSS N l=0.186441u w=1.062u 
.ENDS oai21d1

.SUBCKT oai21d2 ZN  A B1 B2 VDD VSS
MM12 3 2 VDD VDD P l=0.185097u w=1.342u 
MM11 VDD 3 ZN VDD P l=0.184554u w=1.502u 
MM10 VDD 3 ZN VDD P l=0.184861u w=1.506u 
MM9 VDD A 2 VDD P l=0.185213u w=1.312u 
MM8 10 B1 2 VDD P l=0.18u w=1.31u 
MM7 10 B2 VDD VDD P l=0.18u w=1.31u 
MM6 VSS 2 3 VSS N l=0.186381u w=1.072u 
MM5 VSS 3 ZN VSS N l=0.187276u w=1.006u 
MM4 VSS 3 ZN VSS N l=0.186826u w=1.002u 
MM3 2 A 9 VSS N l=0.18u w=1.09u 
MM2 VSS B1 9 VSS N l=0.186441u w=1.062u 
MM1 9 B2 VSS VSS N l=0.186441u w=1.062u 
.ENDS oai21d2

.SUBCKT oai21d4 ZN  A B1 B2 VDD VSS
MM14 VDD 2 3 VDD P l=0.184985u w=1.372u 
MM13 ZN 3 VDD VDD P l=0.183881u w=2.01u 
MM12 ZN 3 VDD VDD P l=0.18516u w=2.035u 
MM11 VDD 3 ZN VDD P l=0.18u w=1.94u 
MM10 VDD A 2 VDD P l=0.185213u w=1.312u 
MM9 10 B1 2 VDD P l=0.18u w=1.31u 
MM8 10 B2 VDD VDD P l=0.18u w=1.31u 
MM7 VSS 2 3 VSS N l=0.186867u w=1.066u 
MM6 ZN 3 VSS VSS N l=0.188286u w=1.383u 
MM5 VSS 3 ZN VSS N l=0.185097u w=1.342u 
MM4 ZN 3 VSS VSS N l=0.18u w=1.28u 
MM3 2 A 9 VSS N l=0.18u w=1.09u 
MM2 VSS B1 9 VSS N l=0.186441u w=1.062u 
MM1 9 B2 VSS VSS N l=0.186441u w=1.062u 
.ENDS oai21d4

.SUBCKT oai221d1 ZN  A B1 B2 C1 C2 VDD VSS
MM10 11 B2 VDD VDD P l=0.18u w=1.38u 
MM9 11 B1 ZN VDD P l=0.18u w=1.38u 
MM8 ZN C1 12 VDD P l=0.18u w=1.38u 
MM7 VDD C2 12 VDD P l=0.18u w=1.38u 
MM6 ZN A VDD VDD P l=0.18u w=1.23u 
MM4 9 B1 10 VSS N l=0.185135u w=1.332u 
MM5 10 B2 9 VSS N l=0.18607u w=1.206u 
MM3 10 A ZN VSS N l=0.18u w=1.14u 
MM2 9 C1 VSS VSS N l=0.186724u w=1.16u 
MM1 9 C2 VSS VSS N l=0.186724u w=1.16u 
.ENDS oai221d1

.SUBCKT oai221d2 ZN  A B1 B2 C1 C2 VDD VSS
MM15 VDD A 4 VDD P l=0.18u w=1.23u 
MM14 VDD 3 ZN VDD P l=0.184711u w=1.452u 
MM13 VDD 3 ZN VDD P l=0.184711u w=1.452u 
MM12 VDD 4 3 VDD P l=0.185342u w=1.46u 
MM11 13 B2 VDD VDD P l=0.18u w=1.38u 
MM10 13 B1 4 VDD P l=0.18u w=1.38u 
MM9 4 C1 14 VDD P l=0.18u w=1.38u 
MM8 VDD C2 14 VDD P l=0.18u w=1.38u 
MM7 10 A 4 VSS N l=0.18u w=1.14u 
MM6 10 B2 12 VSS N l=0.18607u w=1.206u 
MM5 12 B1 10 VSS N l=0.185135u w=1.332u 
MM4 VSS 3 ZN VSS N l=0.198764u w=1.941u 
MM3 VSS 4 3 VSS N l=0.187709u w=1.074u 
MM2 12 C1 VSS VSS N l=0.186724u w=1.16u 
MM1 12 C2 VSS VSS N l=0.186724u w=1.16u 
.ENDS oai221d2

.SUBCKT oai221d4 ZN  A B1 B2 C1 C2 VDD VSS
MM17 VDD A 3 VDD P l=0.18u w=1.23u 
MM16 4 3 VDD VDD P l=0.185597u w=1.222u 
MM15 VDD 4 ZN VDD P l=0.184667u w=1.774u 
MM14 VDD 4 ZN VDD P l=0.18u w=1.7u 
MM13 VDD 4 ZN VDD P l=0.185817u w=1.805u 
MM12 VDD B2 13 VDD P l=0.18u w=1.38u 
MM11 3 B1 13 VDD P l=0.18u w=1.38u 
MM10 3 C1 14 VDD P l=0.18u w=1.38u 
MM9 VDD C2 14 VDD P l=0.18u w=1.38u 
MM8 12 A 3 VSS N l=0.18u w=1.14u 
MM7 12 B2 11 VSS N l=0.18607u w=1.206u 
MM6 11 B1 12 VSS N l=0.185135u w=1.332u 
MM5 4 3 VSS VSS N l=0.186381u w=1.072u 
MM4 VSS 4 ZN VSS N l=0.19031u w=1.775u 
MM3 VSS 4 ZN VSS N l=0.187889u w=1.734u 
MM2 11 C1 VSS VSS N l=0.186724u w=1.16u 
MM1 11 C2 VSS VSS N l=0.186724u w=1.16u 
.ENDS oai221d4

.SUBCKT oai2222d1 ZN  A1 A2 B1 B2 C1 C2 D1 D2 VDD VSS
MM21 4 3 17 VDD P l=0.18u w=1.46u 
MM22 VDD 2 17 VDD P l=0.18u w=1.46u 
MM20 VDD 4 ZN VDD P l=0.18u w=1.5u 
MM19 VDD A2 18 VDD P l=0.18u w=1.44u 
MM18 18 A1 3 VDD P l=0.18u w=0.98u 
MM17 19 B1 3 VDD P l=0.18u w=1.44u 
MM16 19 B2 VDD VDD P l=0.18u w=1.44u 
MM15 20 C1 2 VDD P l=0.18u w=1.44u 
MM14 VDD C2 20 VDD P l=0.18u w=1.44u 
MM12 21 D1 2 VDD P l=0.18u w=1.46u 
MM13 VDD D2 21 VDD P l=0.18u w=1.46u 
MM11 4 2 VSS VSS N l=0.186042u w=1.132u 
MM10 4 3 VSS VSS N l=0.186042u w=1.132u 
MM9 VSS B1 14 VSS N l=0.187238u w=1.144u 
MM8 VSS B2 14 VSS N l=0.186842u w=1.14u 
MM7 ZN 4 VSS VSS N l=0.186826u w=1.002u 
MM6 3 A2 14 VSS N l=0.18u w=1.08u 
MM5 3 A1 14 VSS N l=0.186387u w=1.146u 
MM4 VSS D2 15 VSS N l=0.186042u w=1.132u 
MM3 VSS D1 15 VSS N l=0.186444u w=1.136u 
MM2 2 C1 15 VSS N l=0.1875u w=1.104u 
MM1 2 C2 15 VSS N l=0.187091u w=1.1u 
.ENDS oai2222d1

.SUBCKT oai2222d2 ZN  A1 A2 B1 B2 C1 C2 D1 D2 VDD VSS
MM23 8 3 17 VDD P l=0.18u w=1.46u 
MM24 VDD 2 17 VDD P l=0.18u w=1.46u 
MM22 18 C1 2 VDD P l=0.18u w=1.44u 
MM21 VDD C2 18 VDD P l=0.18u w=1.44u 
MM19 19 D1 2 VDD P l=0.18u w=1.46u 
MM20 VDD D2 19 VDD P l=0.18u w=1.46u 
MM18 VDD 8 ZN VDD P l=0.18u w=1.5u 
MM17 VDD 8 ZN VDD P l=0.18u w=1.5u 
MM16 VDD A2 20 VDD P l=0.18u w=1.44u 
MM15 20 A1 3 VDD P l=0.18u w=0.98u 
MM14 21 B1 3 VDD P l=0.18u w=1.44u 
MM13 21 B2 VDD VDD P l=0.18u w=1.44u 
MM12 8 2 VSS VSS N l=0.186042u w=1.132u 
MM11 8 3 VSS VSS N l=0.186042u w=1.132u 
MM10 VSS B1 14 VSS N l=0.187238u w=1.144u 
MM9 VSS B2 14 VSS N l=0.186842u w=1.14u 
MM8 VSS D2 15 VSS N l=0.186042u w=1.132u 
MM7 VSS D1 15 VSS N l=0.186444u w=1.136u 
MM6 ZN 8 VSS VSS N l=0.186826u w=1.002u 
MM5 ZN 8 VSS VSS N l=0.186826u w=1.002u 
MM4 3 A2 14 VSS N l=0.18u w=1.08u 
MM3 3 A1 14 VSS N l=0.186387u w=1.146u 
MM2 2 C1 15 VSS N l=0.1875u w=1.104u 
MM1 2 C2 15 VSS N l=0.187091u w=1.1u 
.ENDS oai2222d2

.SUBCKT oai2222d4 ZN  A1 A2 B1 B2 C1 C2 D1 D2 VDD VSS
MM26 ZN 2 VDD VDD P l=0.188173u w=2.063u 
MM25 VDD 2 ZN VDD P l=0.18u w=1.91u 
MM24 VDD 2 ZN VDD P l=0.18592u w=2.017u 
MM23 17 D2 VDD VDD P l=0.18u w=1.21u 
MM22 17 D1 12 VDD P l=0.18u w=1.21u 
MM21 18 C1 12 VDD P l=0.18u w=1.21u 
MM20 VDD C2 18 VDD P l=0.18u w=1.21u 
MM19 VDD A2 19 VDD P l=0.18u w=1.21u 
MM18 11 A1 19 VDD P l=0.18u w=1.21u 
MM17 11 B1 20 VDD P l=0.18u w=1.21u 
MM16 VDD B2 20 VDD P l=0.18u w=1.21u 
MM15 2 11 21 VDD P l=0.18u w=1.21u 
MM14 21 12 VDD VDD P l=0.18u w=1.21u 
MM12 VSS 2 ZN VSS N l=0.185656u w=1.464u 
MM13 ZN 2 VSS VSS N l=0.187175u w=1.154u 
MM11 ZN 2 VSS VSS N l=0.18u w=1.39u 
MM10 VSS D2 16 VSS N l=0.18u w=1.08u 
MM9 VSS D1 16 VSS N l=0.186903u w=1.13u 
MM8 2 11 VSS VSS N l=0.18u w=1.06u 
MM7 VSS 12 2 VSS N l=0.186096u w=1.122u 
MM6 15 B1 VSS VSS N l=0.186096u w=1.122u 
MM5 15 B2 VSS VSS N l=0.186096u w=1.122u 
MM3 11 A1 15 VSS N l=0.18u w=0.9u 
MM4 11 A2 15 VSS N l=0.186387u w=1.146u 
MM2 12 C1 16 VSS N l=0.18u w=1.08u 
MM1 12 C2 16 VSS N l=0.186387u w=1.146u 
.ENDS oai2222d4

.SUBCKT oai222d1 ZN  A1 A2 B1 B2 C1 C2 VDD VSS
MM12 VDD B2 12 VDD P l=0.18u w=1.41u 
MM11 ZN B1 12 VDD P l=0.18u w=1.41u 
MM10 ZN C1 13 VDD P l=0.184647u w=1.472u 
MM9 VDD C2 13 VDD P l=0.18527u w=1.48u 
MM8 ZN A1 14 VDD P l=0.188486u w=1.407u 
MM7 VDD A2 14 VDD P l=0.188486u w=1.407u 
MM6 10 B2 11 VSS N l=0.1865u w=1.2u 
MM4 ZN A2 11 VSS N l=0.18u w=1.13u 
MM5 ZN A1 11 VSS N l=0.1865u w=1.2u 
MM3 10 B1 11 VSS N l=0.18u w=1.13u 
MM2 VSS C1 10 VSS N l=0.18u w=1.13u 
MM1 VSS C2 10 VSS N l=0.1865u w=1.2u 
.ENDS oai222d1

.SUBCKT oai222d2 ZN  A1 A2 B1 B2 C1 C2 VDD VSS
MM18 VDD A2 14 VDD P l=0.188486u w=1.407u 
MM17 5 A1 14 VDD P l=0.188486u w=1.407u 
MM16 VDD 4 ZN VDD P l=0.184554u w=1.502u 
MM15 ZN 4 VDD VDD P l=0.184554u w=1.502u 
MM14 4 5 VDD VDD P l=0.186446u w=1.21u 
MM13 VDD B2 15 VDD P l=0.18u w=1.41u 
MM12 5 B1 15 VDD P l=0.18u w=1.41u 
MM11 5 C1 16 VDD P l=0.184647u w=1.472u 
MM10 VDD C2 16 VDD P l=0.18527u w=1.48u 
MM9 5 A2 11 VSS N l=0.18u w=1.13u 
MM7 13 B2 11 VSS N l=0.1865u w=1.2u 
MM8 5 A1 11 VSS N l=0.1865u w=1.2u 
MM6 13 B1 11 VSS N l=0.18u w=1.13u 
MM5 ZN 4 VSS VSS N l=0.186826u w=1.002u 
MM4 ZN 4 VSS VSS N l=0.186826u w=1.002u 
MM3 4 5 VSS VSS N l=0.186381u w=1.072u 
MM2 VSS C1 13 VSS N l=0.18u w=1.13u 
MM1 VSS C2 13 VSS N l=0.1865u w=1.2u 
.ENDS oai222d2

.SUBCKT oai222d4 ZN  A1 A2 B1 B2 C1 C2 VDD VSS
MM19 4 A1 14 VDD P l=0.188486u w=1.407u 
MM18 VDD A2 14 VDD P l=0.188486u w=1.407u 
MM17 5 4 VDD VDD P l=0.18u w=1.44u 
MM16 ZN 5 VDD VDD P l=0.184845u w=1.808u 
MM15 VDD 5 ZN VDD P l=0.18u w=1.73u 
MM14 ZN 5 VDD VDD P l=0.18459u w=1.804u 
MM13 VDD B2 15 VDD P l=0.18u w=1.41u 
MM12 4 B1 15 VDD P l=0.18u w=1.41u 
MM11 4 C1 16 VDD P l=0.184647u w=1.472u 
MM10 VDD C2 16 VDD P l=0.18527u w=1.48u 
MM9 4 A1 11 VSS N l=0.1865u w=1.2u 
MM8 4 A2 11 VSS N l=0.18u w=1.13u 
MM7 13 B2 11 VSS N l=0.1865u w=1.2u 
MM6 13 B1 11 VSS N l=0.18u w=1.13u 
MM5 5 4 VSS VSS N l=0.187222u w=1.08u 
MM4 VSS 5 ZN VSS N l=0.190556u w=1.779u 
MM3 ZN 5 VSS VSS N l=0.190556u w=1.779u 
MM2 VSS C1 13 VSS N l=0.18u w=1.13u 
MM1 VSS C2 13 VSS N l=0.1865u w=1.2u 
.ENDS oai222d4

.SUBCKT oai22d1 ZN  A1 A2 B1 B2 VDD VSS
MM8 VDD A2 9 VDD P l=0.18u w=1.38u 
MM7 ZN A1 9 VDD P l=0.18u w=1.38u 
MM6 10 B1 ZN VDD P l=0.18u w=1.38u 
MM5 VDD B2 10 VDD P l=0.18u w=1.38u 
MM4 8 A2 ZN VSS N l=0.185787u w=1.182u 
MM3 8 A1 ZN VSS N l=0.185787u w=1.182u 
MM2 8 B1 VSS VSS N l=0.18u w=1.12u 
MM1 8 B2 VSS VSS N l=0.186555u w=1.19u 
.ENDS oai22d1

.SUBCKT oai22d2 ZN  A1 A2 B1 B2 VDD VSS
MM14 VDD A2 11 VDD P l=0.18u w=1.38u 
MM13 6 A1 11 VDD P l=0.18u w=1.38u 
MM12 12 B1 6 VDD P l=0.18u w=1.38u 
MM11 VDD B2 12 VDD P l=0.18u w=1.38u 
MM10 7 6 VDD VDD P l=0.185097u w=1.342u 
MM9 ZN 7 VDD VDD P l=0.184554u w=1.502u 
MM8 VDD 7 ZN VDD P l=0.184861u w=1.506u 
MM7 9 A2 6 VSS N l=0.185787u w=1.182u 
MM6 9 A1 6 VSS N l=0.185787u w=1.182u 
MM5 9 B1 VSS VSS N l=0.18u w=1.12u 
MM4 9 B2 VSS VSS N l=0.186555u w=1.19u 
MM3 VSS 6 7 VSS N l=0.186381u w=1.072u 
MM2 ZN 7 VSS VSS N l=0.187276u w=1.006u 
MM1 VSS 7 ZN VSS N l=0.186826u w=1.002u 
.ENDS oai22d2

.SUBCKT oai22d4 ZN  A1 A2 B1 B2 VDD VSS
MM16 3 2 VDD VDD P l=0.184985u w=1.372u 
MM15 VDD 3 ZN VDD P l=0.183881u w=2.01u 
MM14 ZN 3 VDD VDD P l=0.18516u w=2.035u 
MM13 ZN 3 VDD VDD P l=0.18u w=1.94u 
MM12 VDD A2 11 VDD P l=0.18u w=1.38u 
MM11 2 A1 11 VDD P l=0.18u w=1.38u 
MM10 12 B1 2 VDD P l=0.18u w=1.38u 
MM9 VDD B2 12 VDD P l=0.18u w=1.38u 
MM8 VSS 2 3 VSS N l=0.186867u w=1.066u 
MM7 ZN 3 VSS VSS N l=0.188286u w=1.383u 
MM6 VSS 3 ZN VSS N l=0.185097u w=1.342u 
MM5 VSS 3 ZN VSS N l=0.18u w=1.28u 
MM4 10 A2 2 VSS N l=0.185787u w=1.182u 
MM3 10 A1 2 VSS N l=0.185787u w=1.182u 
MM2 10 B1 VSS VSS N l=0.18u w=1.12u 
MM1 10 B2 VSS VSS N l=0.186555u w=1.19u 
.ENDS oai22d4

.SUBCKT oai311d1 ZN  A B C1 C2 C3 VDD VSS
MM10 12 C1 ZN VDD P l=0.18u w=1.97u 
MM7 VDD B ZN VDD P l=0.186441u w=1.062u 
MM9 11 C3 VDD VDD P l=0.18u w=1.97u 
MM8 11 C2 12 VDD P l=0.18u w=1.97u 
MM6 VDD A ZN VDD P l=0.186441u w=1.062u 
MM4 VSS C3 8 VSS N l=0.185836u w=1.172u 
MM3 VSS C2 8 VSS N l=0.185836u w=1.172u 
MM5 VSS C1 8 VSS N l=0.185836u w=1.172u 
MM2 10 B 8 VSS N l=0.18u w=0.97u 
MM1 ZN A 10 VSS N l=0.18u w=0.97u 
.ENDS oai311d1

.SUBCKT oai311d2 ZN  A B C1 C2 C3 VDD VSS
MM14 VDD A 7 VDD P l=0.186441u w=1.062u 
MM16 13 C3 VDD VDD P l=0.18u w=1.97u 
MM13 13 C2 14 VDD P l=0.18u w=1.97u 
MM15 VDD B 7 VDD P l=0.186441u w=1.062u 
MM12 14 C1 7 VDD P l=0.18u w=1.97u 
MM11 VDD 7 8 VDD P l=0.185597u w=1.222u 
MM10 VDD 8 ZN VDD P l=0.184554u w=1.502u 
MM9 VDD 8 ZN VDD P l=0.184554u w=1.502u 
MM7 12 B 11 VSS N l=0.18u w=0.97u 
MM4 VSS C1 11 VSS N l=0.185836u w=1.172u 
MM6 7 A 12 VSS N l=0.18u w=0.97u 
MM8 VSS C3 11 VSS N l=0.185836u w=1.172u 
MM5 VSS C2 11 VSS N l=0.185836u w=1.172u 
MM3 VSS 7 8 VSS N l=0.186381u w=1.072u 
MM2 VSS 8 ZN VSS N l=0.186826u w=1.002u 
MM1 VSS 8 ZN VSS N l=0.186826u w=1.002u 
.ENDS oai311d2

.SUBCKT oai311d4 ZN  A B C1 C2 C3 VDD VSS
MM16 VDD A 7 VDD P l=0.186441u w=1.062u 
MM18 13 C3 VDD VDD P l=0.18u w=1.97u 
MM15 13 C2 14 VDD P l=0.18u w=1.97u 
MM17 VDD B 7 VDD P l=0.186441u w=1.062u 
MM14 14 C1 7 VDD P l=0.18u w=1.97u 
MM13 VDD 7 8 VDD P l=0.185597u w=1.222u 
MM11 ZN 8 VDD VDD P l=0.183417u w=2.002u 
MM12 VDD 8 ZN VDD P l=0.183417u w=2.002u 
MM10 VDD 8 ZN VDD P l=0.183417u w=2.002u 
MM8 12 B 11 VSS N l=0.18u w=0.97u 
MM5 VSS C1 11 VSS N l=0.185836u w=1.172u 
MM7 7 A 12 VSS N l=0.18u w=0.97u 
MM9 VSS C3 11 VSS N l=0.185836u w=1.172u 
MM6 VSS C2 11 VSS N l=0.185836u w=1.172u 
MM4 8 7 VSS VSS N l=0.186381u w=1.072u 
MM3 VSS 8 ZN VSS N l=0.185174u w=1.322u 
MM2 VSS 8 ZN VSS N l=0.185174u w=1.322u 
MM1 VSS 8 ZN VSS N l=0.185059u w=1.352u 
.ENDS oai311d4

.SUBCKT oai31d1 ZN  A B1 B2 B3 VDD VSS
MM8 10 B2 9 VDD P l=0.18u w=1.71u 
MM7 VDD B3 9 VDD P l=0.18u w=1.71u 
MM6 ZN A VDD VDD P l=0.18u w=0.97u 
MM5 ZN B1 10 VDD P l=0.18u w=1.71u 
MM4 VSS B2 7 VSS N l=0.187066u w=1.036u 
MM3 VSS B3 7 VSS N l=0.1878u w=1u 
MM2 7 A ZN VSS N l=0.18u w=0.9u 
MM1 VSS B1 7 VSS N l=0.18u w=0.9u 
.ENDS oai31d1

.SUBCKT oai31d2 ZN  A B1 B2 B3 VDD VSS
MM14 3 2 VDD VDD P l=0.185097u w=1.342u 
MM13 ZN 3 VDD VDD P l=0.184554u w=1.502u 
MM12 VDD 3 ZN VDD P l=0.184861u w=1.506u 
MM11 VDD B3 11 VDD P l=0.18u w=1.71u 
MM9 12 B2 11 VDD P l=0.18u w=1.71u 
MM10 2 A VDD VDD P l=0.18u w=1.34u 
MM8 2 B1 12 VDD P l=0.18u w=1.71u 
MM6 2 A 10 VSS N l=0.186441u w=1.062u 
MM7 10 B3 VSS VSS N l=0.18u w=1.04u 
MM5 VSS B2 10 VSS N l=0.186502u w=1.052u 
MM4 VSS B1 10 VSS N l=0.18u w=1u 
MM3 VSS 2 3 VSS N l=0.186381u w=1.072u 
MM2 VSS 3 ZN VSS N l=0.187276u w=1.006u 
MM1 VSS 3 ZN VSS N l=0.186826u w=1.002u 
.ENDS oai31d2

.SUBCKT oai31d4 ZN  A B1 B2 B3 VDD VSS
MM16 3 2 VDD VDD P l=0.184985u w=1.372u 
MM15 VDD 3 ZN VDD P l=0.183881u w=2.01u 
MM14 ZN 3 VDD VDD P l=0.18516u w=2.035u 
MM13 ZN 3 VDD VDD P l=0.18u w=1.94u 
MM11 11 B3 VDD VDD P l=0.18u w=1.71u 
MM10 11 B2 12 VDD P l=0.18u w=1.71u 
MM12 2 A VDD VDD P l=0.18u w=0.97u 
MM9 2 B1 12 VDD P l=0.18u w=1.71u 
MM8 VSS 2 3 VSS N l=0.186322u w=1.082u 
MM7 VSS 3 ZN VSS N l=0.188286u w=1.383u 
MM6 VSS 3 ZN VSS N l=0.185097u w=1.342u 
MM5 ZN 3 VSS VSS N l=0.18u w=1.28u 
MM4 2 A 10 VSS N l=0.186502u w=1.052u 
MM3 10 B3 VSS VSS N l=0.18u w=1.04u 
MM2 VSS B2 10 VSS N l=0.186932u w=1.056u 
MM1 VSS B1 10 VSS N l=0.18u w=0.99u 
.ENDS oai31d4

.SUBCKT oai321d1 ZN  A B1 B2 C1 C2 C3 VDD VSS
MM11 ZN A VDD VDD P l=0.187528u w=1.331u 
MM12 ZN B1 12 VDD P l=0.18u w=1.24u 
MM10 12 B2 VDD VDD P l=0.18u w=1.24u 
MM9 13 C3 VDD VDD P l=0.18u w=1.24u 
MM7 13 C2 14 VDD P l=0.18u w=1.24u 
MM8 ZN C1 14 VDD P l=0.18u w=1.24u 
MM6 10 B1 11 VSS N l=0.184679u w=1.462u 
MM5 11 A ZN VSS N l=0.186502u w=1.052u 
MM4 11 B2 10 VSS N l=0.18u w=0.9u 
MM2 10 C1 VSS VSS N l=0.186387u w=1.146u 
MM3 VSS C3 10 VSS N l=0.186783u w=1.15u 
MM1 VSS C2 10 VSS N l=0.18u w=1.08u 
.ENDS oai321d1

.SUBCKT oai321d2 ZN  A B1 B2 C1 C2 C3 VDD VSS
MM17 8 A VDD VDD P l=0.187528u w=1.331u 
MM16 14 C3 VDD VDD P l=0.18u w=1.24u 
MM13 14 C2 16 VDD P l=0.18u w=1.24u 
MM18 15 B2 VDD VDD P l=0.18u w=1.24u 
MM15 8 B1 15 VDD P l=0.18u w=1.24u 
MM14 8 C1 16 VDD P l=0.18u w=1.24u 
MM12 VDD 8 9 VDD P l=0.185597u w=1.222u 
MM11 VDD 9 ZN VDD P l=0.184554u w=1.502u 
MM10 VDD 9 ZN VDD P l=0.184554u w=1.502u 
MM9 11 B2 13 VSS N l=0.18u w=0.9u 
MM7 13 B1 11 VSS N l=0.184679u w=1.462u 
MM8 11 A 8 VSS N l=0.186502u w=1.052u 
MM6 VSS 8 9 VSS N l=0.186381u w=1.072u 
MM5 ZN 9 VSS VSS N l=0.186826u w=1.002u 
MM4 ZN 9 VSS VSS N l=0.186826u w=1.002u 
MM2 13 C1 VSS VSS N l=0.186387u w=1.146u 
MM3 VSS C3 13 VSS N l=0.186783u w=1.15u 
MM1 VSS C2 13 VSS N l=0.18u w=1.08u 
.ENDS oai321d2

.SUBCKT oai321d4 ZN  A B1 B2 C1 C2 C3 VDD VSS
MM20 8 A VDD VDD P l=0.187528u w=1.331u 
MM19 14 C3 VDD VDD P l=0.18u w=1.24u 
MM15 14 C2 16 VDD P l=0.18u w=1.24u 
MM18 15 B2 VDD VDD P l=0.18u w=1.24u 
MM17 8 B1 15 VDD P l=0.18u w=1.24u 
MM16 8 C1 16 VDD P l=0.18u w=1.24u 
MM14 VDD 8 9 VDD P l=0.185597u w=1.222u 
MM12 VDD 9 ZN VDD P l=0.183417u w=2.002u 
MM13 VDD 9 ZN VDD P l=0.183417u w=2.002u 
MM11 ZN 9 VDD VDD P l=0.183417u w=2.002u 
MM10 13 A 8 VSS N l=0.186502u w=1.052u 
MM9 13 B2 12 VSS N l=0.18u w=0.9u 
MM8 12 B1 13 VSS N l=0.184679u w=1.462u 
MM7 VSS 8 9 VSS N l=0.186381u w=1.072u 
MM6 VSS 9 ZN VSS N l=0.185135u w=1.332u 
MM5 ZN 9 VSS VSS N l=0.185135u w=1.332u 
MM4 VSS 9 ZN VSS N l=0.185135u w=1.332u 
MM2 12 C1 VSS VSS N l=0.186387u w=1.146u 
MM3 VSS C3 12 VSS N l=0.186783u w=1.15u 
MM1 VSS C2 12 VSS N l=0.18u w=1.08u 
.ENDS oai321d4

.SUBCKT oai322d1 ZN  A1 A2 B1 B2 C1 C2 C3 VDD VSS
MM14 13 C3 VDD VDD P l=0.18u w=1.35u 
MM13 13 C2 14 VDD P l=0.18u w=1.35u 
MM12 ZN C1 14 VDD P l=0.18u w=1.35u 
MM9 ZN B1 16 VDD P l=0.18u w=1.2u 
MM11 VDD A2 15 VDD P l=0.18u w=1.11u 
MM10 15 A1 ZN VDD P l=0.18u w=1.11u 
MM8 VDD B2 16 VDD P l=0.18u w=1.2u 
MM7 ZN A2 12 VSS N l=0.18u w=1.09u 
MM6 ZN A1 12 VSS N l=0.186724u w=1.16u 
MM5 12 B1 11 VSS N l=0.18u w=1.38u 
MM4 12 B2 11 VSS N l=0.184743u w=1.442u 
MM3 VSS C3 11 VSS N l=0.186555u w=1.19u 
MM2 VSS C2 11 VSS N l=0.18u w=1.12u 
MM1 VSS C1 11 VSS N l=0.190445u w=1.235u 
.ENDS oai322d1

.SUBCKT oai322d2 ZN  A1 A2 B1 B2 C1 C2 C3 VDD VSS
MM18 4 C1 15 VDD P l=0.18u w=1.35u 
MM13 4 B1 18 VDD P l=0.18u w=1.2u 
MM19 15 C2 16 VDD P l=0.18u w=1.35u 
MM17 10 4 VDD VDD P l=0.18u w=1.35u 
MM16 16 C3 VDD VDD P l=0.18u w=1.35u 
MM15 VDD A2 17 VDD P l=0.18u w=1.15u 
MM14 17 A1 4 VDD P l=0.18u w=1.15u 
MM12 VDD B2 18 VDD P l=0.18u w=1.2u 
MM11 VDD 10 ZN VDD P l=0.18u w=1.38u 
MM10 VDD 10 ZN VDD P l=0.18u w=1.38u 
MM8 VSS C1 12 VSS N l=0.190445u w=1.235u 
MM7 10 4 VSS VSS N l=0.18u w=1.24u 
MM9 VSS C2 12 VSS N l=0.18u w=1.12u 
MM6 VSS C3 12 VSS N l=0.186935u w=1.194u 
MM5 ZN 10 VSS VSS N l=0.193916u w=1.841u 
MM4 4 A2 14 VSS N l=0.18u w=1.09u 
MM3 4 A1 14 VSS N l=0.186724u w=1.16u 
MM2 14 B1 12 VSS N l=0.18u w=1.38u 
MM1 14 B2 12 VSS N l=0.184743u w=1.442u 
.ENDS oai322d2

.SUBCKT oai322d4 ZN  A1 A2 B1 B2 C1 C2 C3 VDD VSS
MM20 10 3 VDD VDD P l=0.18u w=1.35u 
MM21 18 C2 15 VDD P l=0.18u w=1.35u 
MM19 15 C3 VDD VDD P l=0.18u w=1.35u 
MM18 VDD A2 16 VDD P l=0.18u w=1.15u 
MM17 16 A1 3 VDD P l=0.18u w=1.15u 
MM16 3 B1 17 VDD P l=0.18u w=1.2u 
MM14 18 C1 3 VDD P l=0.18u w=1.35u 
MM15 VDD B2 17 VDD P l=0.18u w=1.2u 
MM13 VDD 10 ZN VDD P l=0.189649u w=1.797u 
MM12 VDD 10 ZN VDD P l=0.18u w=1.64u 
MM11 VDD 10 ZN VDD P l=0.186314u w=1.739u 
MM9 10 3 VSS VSS N l=0.18u w=1.24u 
MM10 VSS C2 12 VSS N l=0.18u w=1.12u 
MM8 VSS C3 12 VSS N l=0.186935u w=1.194u 
MM7 VSS C1 12 VSS N l=0.190445u w=1.235u 
MM6 ZN 10 VSS VSS N l=0.187889u w=1.734u 
MM5 ZN 10 VSS VSS N l=0.187217u w=1.721u 
MM4 3 A2 14 VSS N l=0.18u w=1.09u 
MM3 3 A1 14 VSS N l=0.186724u w=1.16u 
MM2 14 B1 12 VSS N l=0.18u w=1.38u 
MM1 14 B2 12 VSS N l=0.184743u w=1.442u 
.ENDS oai322d4

.SUBCKT oaim211d1 ZN  A B C1 C2 VDD VSS
MM9 ZN A VDD VDD P l=0.18u w=1.2u 
MM10 VDD B ZN VDD P l=0.185738u w=1.192u 
MM8 VDD 4 ZN VDD P l=0.185738u w=1.192u 
MM7 4 C2 VDD VDD P l=0.18u w=1.13u 
MM6 4 C1 VDD VDD P l=0.187252u w=1.208u 
MM4 ZN A 9 VSS N l=0.18u w=1.27u 
MM5 10 B 9 VSS N l=0.18u w=1.27u 
MM3 VSS 4 10 VSS N l=0.18u w=1.27u 
MM2 VSS C2 11 VSS N l=0.18u w=0.9u 
MM1 11 C1 4 VSS N l=0.18u w=0.9u 
.ENDS oaim211d1

.SUBCKT oaim211d2 ZN  A B C1 C2 VDD VSS
MM16 7 A VDD VDD P l=0.18u w=1.2u 
MM15 VDD B 7 VDD P l=0.185738u w=1.192u 
MM14 VDD 4 7 VDD P l=0.185738u w=1.192u 
MM13 4 C2 VDD VDD P l=0.18u w=1.13u 
MM12 4 C1 VDD VDD P l=0.187252u w=1.208u 
MM11 VDD 7 8 VDD P l=0.185597u w=1.222u 
MM10 ZN 8 VDD VDD P l=0.184436u w=1.542u 
MM9 VDD 8 ZN VDD P l=0.18u w=1.54u 
MM8 7 A 11 VSS N l=0.18u w=1.27u 
MM7 12 B 11 VSS N l=0.18u w=1.27u 
MM6 VSS 4 12 VSS N l=0.18u w=1.27u 
MM5 VSS C2 13 VSS N l=0.18u w=0.9u 
MM4 13 C1 4 VSS N l=0.18u w=0.9u 
MM3 8 7 VSS VSS N l=0.186381u w=1.072u 
MM2 VSS 8 ZN VSS N l=0.186628u w=1.032u 
MM1 ZN 8 VSS VSS N l=0.186628u w=1.032u 
.ENDS oaim211d2

.SUBCKT oaim211d4 ZN  A B C1 C2 VDD VSS
MM17 VDD B 7 VDD P l=0.185738u w=1.192u 
MM16 VDD 3 7 VDD P l=0.185738u w=1.192u 
MM15 3 C2 VDD VDD P l=0.18u w=1.13u 
MM14 3 C1 VDD VDD P l=0.187252u w=1.208u 
MM13 7 A VDD VDD P l=0.18u w=1.2u 
MM12 VDD 7 8 VDD P l=0.18u w=1.21u 
MM11 ZN 8 VDD VDD P l=0.183713u w=1.842u 
MM10 ZN 8 VDD VDD P l=0.183713u w=1.842u 
MM9 ZN 8 VDD VDD P l=0.18u w=1.78u 
MM8 11 B 13 VSS N l=0.18u w=1.27u 
MM7 VSS 3 11 VSS N l=0.18u w=1.27u 
MM6 VSS C2 12 VSS N l=0.18u w=0.9u 
MM5 12 C1 3 VSS N l=0.18u w=0.9u 
MM4 7 A 13 VSS N l=0.18u w=1.27u 
MM3 8 7 VSS VSS N l=0.186381u w=1.072u 
MM2 VSS 8 ZN VSS N l=0.194726u w=1.858u 
MM1 VSS 8 ZN VSS N l=0.19031u w=1.775u 
.ENDS oaim211d4

.SUBCKT oaim21d1 ZN  A B1 B2 VDD VSS
MM8 VDD A ZN VDD P l=0.185989u w=1.142u 
MM7 VDD 3 ZN VDD P l=0.185989u w=1.142u 
MM6 VDD B2 3 VDD P l=0.186387u w=1.146u 
MM5 VDD B1 3 VDD P l=0.18u w=1.08u 
MM4 8 A ZN VSS N l=0.18u w=0.98u 
MM3 8 3 VSS VSS N l=0.18u w=0.98u 
MM2 9 B2 VSS VSS N l=0.18u w=0.98u 
MM1 3 B1 9 VSS N l=0.18u w=0.98u 
.ENDS oaim21d1

.SUBCKT oaim21d2 ZN  A B1 B2 VDD VSS
MM14 VDD A 6 VDD P l=0.185989u w=1.142u 
MM13 VDD 3 6 VDD P l=0.185989u w=1.142u 
MM12 VDD B2 3 VDD P l=0.186387u w=1.146u 
MM11 VDD B1 3 VDD P l=0.18u w=1.08u 
MM10 7 6 VDD VDD P l=0.185597u w=1.222u 
MM9 VDD 7 ZN VDD P l=0.184554u w=1.502u 
MM8 ZN 7 VDD VDD P l=0.184554u w=1.502u 
MM7 10 A 6 VSS N l=0.18u w=0.98u 
MM6 10 3 VSS VSS N l=0.18u w=0.98u 
MM5 11 B2 VSS VSS N l=0.18u w=0.98u 
MM4 3 B1 11 VSS N l=0.18u w=0.98u 
MM3 VSS 6 7 VSS N l=0.186381u w=1.072u 
MM2 VSS 7 ZN VSS N l=0.186826u w=1.002u 
MM1 VSS 7 ZN VSS N l=0.186826u w=1.002u 
.ENDS oaim21d2

.SUBCKT oaim21d4 ZN  A B1 B2 VDD VSS
MM16 3 2 VDD VDD P l=0.185597u w=1.222u 
MM14 VDD 3 ZN VDD P l=0.183417u w=2.002u 
MM15 ZN 3 VDD VDD P l=0.183417u w=2.002u 
MM13 ZN 3 VDD VDD P l=0.183417u w=2.002u 
MM12 VDD A 2 VDD P l=0.185989u w=1.142u 
MM11 VDD 5 2 VDD P l=0.185989u w=1.142u 
MM10 VDD B2 5 VDD P l=0.186387u w=1.146u 
MM9 VDD B1 5 VDD P l=0.18u w=1.08u 
MM8 VSS 2 3 VSS N l=0.186381u w=1.072u 
MM7 ZN 3 VSS VSS N l=0.185135u w=1.332u 
MM6 VSS 3 ZN VSS N l=0.185135u w=1.332u 
MM5 VSS 3 ZN VSS N l=0.185135u w=1.332u 
MM4 10 A 2 VSS N l=0.18u w=0.98u 
MM3 10 5 VSS VSS N l=0.18u w=0.98u 
MM2 11 B2 VSS VSS N l=0.18u w=0.98u 
MM1 5 B1 11 VSS N l=0.18u w=0.98u 
.ENDS oaim21d4

.SUBCKT oaim22d1 ZN  A1 A2 B1 B2 VDD VSS
MM10 VDD 2 ZN VDD P l=0.18u w=1.18u 
MM8 11 A1 ZN VDD P l=0.18u w=1.51u 
MM9 11 A2 VDD VDD P l=0.18u w=1.51u 
MM7 VDD B2 2 VDD P l=0.185507u w=1.242u 
MM6 VDD B1 2 VDD P l=0.185507u w=1.242u 
MM5 VSS 2 9 VSS N l=0.18u w=1.15u 
MM3 9 A1 ZN VSS N l=0.186501u w=1.126u 
MM4 9 A2 ZN VSS N l=0.18729u w=1.07u 
MM2 VSS B2 10 VSS N l=0.18u w=0.9u 
MM1 10 B1 2 VSS N l=0.18u w=0.9u 
.ENDS oaim22d1

.SUBCKT oaim22d2 ZN  A1 A2 B1 B2 VDD VSS
MM14 VDD B2 3 VDD P l=0.185174u w=1.322u 
MM13 VDD B1 3 VDD P l=0.185174u w=1.322u 
MM15 VDD 3 7 VDD P l=0.18u w=1.26u 
MM12 13 A1 7 VDD P l=0.18u w=1.51u 
MM16 VDD A2 13 VDD P l=0.18u w=1.51u 
MM11 VDD 7 8 VDD P l=0.185335u w=1.282u 
MM10 ZN 8 VDD VDD P l=0.184554u w=1.502u 
MM9 VDD 8 ZN VDD P l=0.184554u w=1.502u 
MM8 10 A2 7 VSS N l=0.187156u w=1.09u 
MM7 10 3 VSS VSS N l=0.18u w=1.15u 
MM4 10 A1 7 VSS N l=0.186444u w=1.136u 
MM6 VSS B2 12 VSS N l=0.18u w=0.9u 
MM5 12 B1 3 VSS N l=0.18u w=0.9u 
MM3 VSS 7 8 VSS N l=0.186441u w=1.062u 
MM2 VSS 8 ZN VSS N l=0.186826u w=1.002u 
MM1 ZN 8 VSS VSS N l=0.186826u w=1.002u 
.ENDS oaim22d2

.SUBCKT oaim22d4 ZN  A1 A2 B1 B2 VDD VSS
MM15 VDD B2 3 VDD P l=0.185174u w=1.322u 
MM14 VDD B1 3 VDD P l=0.185174u w=1.322u 
MM16 VDD 3 7 VDD P l=0.18u w=1.26u 
MM13 13 A1 7 VDD P l=0.18u w=1.51u 
MM17 VDD A2 13 VDD P l=0.18u w=1.51u 
MM12 VDD 7 8 VDD P l=0.185335u w=1.282u 
MM11 ZN 8 VDD VDD P l=0.183615u w=1.892u 
MM10 ZN 8 VDD VDD P l=0.183615u w=1.892u 
MM9 VDD 8 ZN VDD P l=0.183615u w=1.892u 
MM8 10 A2 7 VSS N l=0.186264u w=1.092u 
MM7 10 3 VSS VSS N l=0.18u w=1.15u 
MM4 10 A1 7 VSS N l=0.186444u w=1.136u 
MM6 VSS B2 12 VSS N l=0.18u w=0.9u 
MM5 12 B1 3 VSS N l=0.18u w=0.9u 
MM3 VSS 7 8 VSS N l=0.185022u w=1.362u 
MM2 VSS 8 ZN VSS N l=0.193769u w=2.022u 
MM1 VSS 8 ZN VSS N l=0.190556u w=1.779u 
.ENDS oaim22d4

.SUBCKT oaim2m11d1 ZN  A B C1 C2 VDD VSS
MM11 ZN A VDD VDD P l=0.185836u w=1.172u 
MM10 6 C2 VDD VDD P l=0.187302u w=1.134u 
MM9 6 C1 VDD VDD P l=0.186501u w=1.126u 
MM12 ZN 2 VDD VDD P l=0.187374u w=1.188u 
MM8 ZN 6 VDD VDD P l=0.18u w=1.11u 
MM7 VDD B 2 VDD P l=0.18u w=0.58u 
MM5 10 A ZN VSS N l=0.18u w=0.96u 
MM6 12 2 10 VSS N l=0.18u w=0.96u 
MM4 11 C2 VSS VSS N l=0.18u w=0.96u 
MM3 11 C1 6 VSS N l=0.18u w=0.96u 
MM2 VSS 6 12 VSS N l=0.18u w=0.96u 
MM1 VSS B 2 VSS N l=0.18u w=0.48u 
.ENDS oaim2m11d1

.SUBCKT oaim2m11d2 ZN  A B C1 C2 VDD VSS
MM18 5 B VDD VDD P l=0.18u w=0.58u 
MM17 4 3 VDD VDD P l=0.185597u w=1.222u 
MM16 VDD 4 ZN VDD P l=0.184554u w=1.502u 
MM15 VDD 4 ZN VDD P l=0.184554u w=1.502u 
MM13 9 C2 VDD VDD P l=0.187302u w=1.134u 
MM12 9 C1 VDD VDD P l=0.186501u w=1.126u 
MM11 VDD A 3 VDD P l=0.185836u w=1.172u 
MM14 VDD 5 3 VDD P l=0.187374u w=1.188u 
MM10 3 9 VDD VDD P l=0.18u w=1.11u 
MM9 VSS B 5 VSS N l=0.18u w=0.48u 
MM7 VSS C2 12 VSS N l=0.18u w=0.96u 
MM6 12 C1 9 VSS N l=0.18u w=0.96u 
MM5 13 A 3 VSS N l=0.18u w=0.96u 
MM8 14 5 13 VSS N l=0.18u w=0.96u 
MM4 VSS 9 14 VSS N l=0.18u w=0.96u 
MM3 4 3 VSS VSS N l=0.186381u w=1.072u 
MM2 VSS 4 ZN VSS N l=0.186826u w=1.002u 
MM1 VSS 4 ZN VSS N l=0.186826u w=1.002u 
.ENDS oaim2m11d2

.SUBCKT oaim2m11d4 ZN  A B C1 C2 VDD VSS
MM20 3 2 VDD VDD P l=0.18u w=1.22u 
MM18 ZN 3 VDD VDD P l=0.183417u w=2.002u 
MM19 VDD 3 ZN VDD P l=0.183417u w=2.002u 
MM17 VDD 3 ZN VDD P l=0.183417u w=2.002u 
MM16 VDD B 5 VDD P l=0.18u w=0.58u 
MM14 9 C2 VDD VDD P l=0.187302u w=1.134u 
MM13 9 C1 VDD VDD P l=0.186501u w=1.126u 
MM12 VDD A 2 VDD P l=0.185836u w=1.172u 
MM15 VDD 5 2 VDD P l=0.187374u w=1.188u 
MM11 2 9 VDD VDD P l=0.18u w=1.11u 
MM10 3 2 VSS VSS N l=0.186381u w=1.072u 
MM9 VSS 3 ZN VSS N l=0.185135u w=1.332u 
MM8 VSS 3 ZN VSS N l=0.185135u w=1.332u 
MM7 ZN 3 VSS VSS N l=0.185135u w=1.332u 
MM6 5 B VSS VSS N l=0.18u w=0.48u 
MM4 VSS C2 12 VSS N l=0.18u w=0.96u 
MM3 12 C1 9 VSS N l=0.18u w=0.96u 
MM2 13 A 2 VSS N l=0.18u w=0.96u 
MM5 14 5 13 VSS N l=0.18u w=0.96u 
MM1 VSS 9 14 VSS N l=0.18u w=0.96u 
.ENDS oaim2m11d4

.SUBCKT oaim311d1 ZN  A B C1 C2 C3 VDD VSS
MM11 ZN A VDD VDD P l=0.185954u w=1.31u 
MM12 ZN 2 VDD VDD P l=0.18u w=1.24u 
MM10 ZN B VDD VDD P l=0.185954u w=1.31u 
MM9 2 C3 VDD VDD P l=0.185479u w=1.336u 
MM8 2 C2 VDD VDD P l=0.18u w=1.27u 
MM7 2 C1 VDD VDD P l=0.185821u w=1.34u 
MM5 ZN A 10 VSS N l=0.18u w=0.96u 
MM4 11 B 10 VSS N l=0.18u w=0.96u 
MM6 VSS 2 11 VSS N l=0.18u w=0.96u 
MM3 VSS C3 12 VSS N l=0.18u w=0.96u 
MM2 13 C2 12 VSS N l=0.18u w=0.96u 
MM1 13 C1 2 VSS N l=0.18u w=0.96u 
.ENDS oaim311d1

.SUBCKT oaim311d2 ZN  A B C1 C2 C3 VDD VSS
MM18 VDD A 8 VDD P l=0.185954u w=1.31u 
MM16 3 C3 VDD VDD P l=0.185479u w=1.336u 
MM15 3 C2 VDD VDD P l=0.18u w=1.27u 
MM14 3 C1 VDD VDD P l=0.185821u w=1.34u 
MM17 8 3 VDD VDD P l=0.18u w=1.24u 
MM13 8 B VDD VDD P l=0.18u w=1.31u 
MM12 VDD 8 9 VDD P l=0.185097u w=1.342u 
MM11 VDD 9 ZN VDD P l=0.185696u w=1.538u 
MM10 VDD 9 ZN VDD P l=0.18u w=1.46u 
MM9 8 A 14 VSS N l=0.18u w=0.96u 
MM7 VSS C3 12 VSS N l=0.18u w=0.96u 
MM6 13 C2 12 VSS N l=0.18u w=0.96u 
MM5 13 C1 3 VSS N l=0.18u w=0.96u 
MM4 14 B 15 VSS N l=0.18u w=0.96u 
MM8 VSS 3 15 VSS N l=0.18u w=0.96u 
MM3 VSS 8 9 VSS N l=0.186381u w=1.072u 
MM2 VSS 9 ZN VSS N l=0.186502u w=1.052u 
MM1 VSS 9 ZN VSS N l=0.18u w=0.94u 
.ENDS oaim311d2

.SUBCKT oaim311d4 ZN  A B C1 C2 C3 VDD VSS
MM20 VDD A 8 VDD P l=0.185954u w=1.31u 
MM18 3 C3 VDD VDD P l=0.185479u w=1.336u 
MM17 3 C2 VDD VDD P l=0.18u w=1.27u 
MM16 3 C1 VDD VDD P l=0.185821u w=1.34u 
MM19 8 3 VDD VDD P l=0.18u w=1.24u 
MM15 8 B VDD VDD P l=0.18u w=1.31u 
MM14 9 8 VDD VDD P l=0.184985u w=1.372u 
MM13 ZN 9 VDD VDD P l=0.183881u w=2.01u 
MM12 VDD 9 ZN VDD P l=0.184111u w=2.014u 
MM11 VDD 9 ZN VDD P l=0.18u w=1.94u 
MM10 8 A 14 VSS N l=0.18u w=0.96u 
MM8 VSS C3 12 VSS N l=0.18u w=0.96u 
MM7 13 C2 12 VSS N l=0.18u w=0.96u 
MM6 13 C1 3 VSS N l=0.18u w=0.96u 
MM5 14 B 15 VSS N l=0.18u w=0.96u 
MM9 VSS 3 15 VSS N l=0.18u w=0.96u 
MM4 VSS 8 9 VSS N l=0.189991u w=1.099u 
MM2 ZN 9 VSS VSS N l=0.185778u w=1.35u 
MM3 ZN 9 VSS VSS N l=0.185097u w=1.342u 
MM1 ZN 9 VSS VSS N l=0.18u w=1.28u 
.ENDS oaim311d4

.SUBCKT oaim31d1 ZN  A B1 B2 B3 VDD VSS
MM9 ZN A VDD VDD P l=0.184985u w=1.372u 
MM8 ZN 4 VDD VDD P l=0.184985u w=1.372u 
MM7 4 B1 VDD VDD P l=0.185213u w=1.312u 
MM10 VDD B3 4 VDD P l=0.18u w=1.31u 
MM6 VDD B2 4 VDD P l=0.184985u w=1.372u 
MM4 ZN A 9 VSS N l=0.18u w=0.86u 
MM3 VSS 4 9 VSS N l=0.18u w=0.86u 
MM2 11 B1 4 VSS N l=0.18u w=0.81u 
MM5 VSS B3 10 VSS N l=0.18u w=0.81u 
MM1 11 B2 10 VSS N l=0.18u w=0.81u 
.ENDS oaim31d1

.SUBCKT oaim31d2 ZN  A B1 B2 B3 VDD VSS
MM15 6 B1 VDD VDD P l=0.185213u w=1.312u 
MM14 VDD B2 6 VDD P l=0.184985u w=1.372u 
MM13 VDD B3 6 VDD P l=0.18u w=1.31u 
MM16 7 A VDD VDD P l=0.184985u w=1.372u 
MM12 7 6 VDD VDD P l=0.184985u w=1.372u 
MM11 VDD 7 8 VDD P l=0.185097u w=1.342u 
MM10 VDD 8 ZN VDD P l=0.184554u w=1.502u 
MM9 VDD 8 ZN VDD P l=0.184861u w=1.506u 
MM8 7 A 13 VSS N l=0.18u w=0.86u 
MM7 11 B1 6 VSS N l=0.18u w=0.81u 
MM6 11 B2 12 VSS N l=0.18u w=0.81u 
MM5 VSS B3 12 VSS N l=0.18u w=0.81u 
MM4 VSS 6 13 VSS N l=0.18u w=0.86u 
MM3 8 7 VSS VSS N l=0.186381u w=1.072u 
MM2 VSS 8 ZN VSS N l=0.187276u w=1.006u 
MM1 VSS 8 ZN VSS N l=0.186826u w=1.002u 
.ENDS oaim31d2

.SUBCKT oaim31d4 ZN  A B1 B2 B3 VDD VSS
MM17 6 B1 VDD VDD P l=0.185213u w=1.312u 
MM16 VDD B2 6 VDD P l=0.184985u w=1.372u 
MM15 VDD B3 6 VDD P l=0.18u w=1.31u 
MM18 7 A VDD VDD P l=0.184985u w=1.372u 
MM14 7 6 VDD VDD P l=0.184985u w=1.372u 
MM13 VDD 7 8 VDD P l=0.184985u w=1.372u 
MM12 VDD 8 ZN VDD P l=0.183881u w=2.01u 
MM11 VDD 8 ZN VDD P l=0.18516u w=2.035u 
MM10 VDD 8 ZN VDD P l=0.18u w=1.94u 
MM9 7 A 13 VSS N l=0.18u w=0.86u 
MM8 11 B1 6 VSS N l=0.18u w=0.81u 
MM7 11 B2 12 VSS N l=0.18u w=0.81u 
MM6 VSS B3 12 VSS N l=0.18u w=0.81u 
MM5 VSS 6 13 VSS N l=0.18u w=0.86u 
MM4 8 7 VSS VSS N l=0.186867u w=1.066u 
MM3 VSS 8 ZN VSS N l=0.188286u w=1.383u 
MM2 ZN 8 VSS VSS N l=0.185097u w=1.342u 
MM1 ZN 8 VSS VSS N l=0.18u w=1.28u 
.ENDS oaim31d4

.SUBCKT oaim3m11d1 ZN  A B C1 C2 C3 VDD VSS
MM13 ZN A VDD VDD P l=0.186207u w=1.102u 
MM14 VDD 2 ZN VDD P l=0.186679u w=1.096u 
MM12 VDD 4 ZN VDD P l=0.18u w=1.03u 
MM11 VDD C2 4 VDD P l=0.18u w=1.08u 
MM10 VDD C3 4 VDD P l=0.18u w=1.15u 
MM9 VDD C1 4 VDD P l=0.18u w=1.15u 
MM8 VDD B 2 VDD P l=0.18u w=0.5u 
MM6 ZN A 11 VSS N l=0.18u w=0.98u 
MM7 11 2 12 VSS N l=0.18u w=0.98u 
MM5 VSS 4 12 VSS N l=0.18u w=0.98u 
MM4 13 C2 14 VSS N l=0.18u w=0.98u 
MM3 13 C3 VSS VSS N l=0.18u w=0.98u 
MM2 4 C1 14 VSS N l=0.18u w=0.98u 
MM1 VSS B 2 VSS N l=0.18u w=0.48u 
.ENDS oaim3m11d1

.SUBCKT oaim3m11d2 ZN  A B C1 C2 C3 VDD VSS
MM20 VDD 2 8 VDD P l=0.186679u w=1.096u 
MM19 VDD 3 8 VDD P l=0.18u w=1.03u 
MM18 8 A VDD VDD P l=0.186207u w=1.102u 
MM17 VDD C2 3 VDD P l=0.18u w=1.08u 
MM16 VDD C3 3 VDD P l=0.18u w=1.15u 
MM15 VDD C1 3 VDD P l=0.18u w=1.15u 
MM14 9 8 VDD VDD P l=0.185097u w=1.342u 
MM13 ZN 9 VDD VDD P l=0.184554u w=1.502u 
MM12 VDD 9 ZN VDD P l=0.184861u w=1.506u 
MM11 VDD B 2 VDD P l=0.18u w=0.5u 
MM10 9 8 VSS VSS N l=0.186381u w=1.072u 
MM9 ZN 9 VSS VSS N l=0.187276u w=1.006u 
MM8 ZN 9 VSS VSS N l=0.186826u w=1.002u 
MM7 14 2 13 VSS N l=0.18u w=0.98u 
MM6 VSS 3 13 VSS N l=0.18u w=0.98u 
MM5 8 A 14 VSS N l=0.18u w=0.98u 
MM4 15 C2 16 VSS N l=0.18u w=0.98u 
MM3 15 C3 VSS VSS N l=0.18u w=0.98u 
MM2 3 C1 16 VSS N l=0.18u w=0.98u 
MM1 VSS B 2 VSS N l=0.18u w=0.48u 
.ENDS oaim3m11d2

.SUBCKT oaim3m11d4 ZN  A B C1 C2 C3 VDD VSS
MM22 3 2 VDD VDD P l=0.184985u w=1.372u 
MM21 VDD 3 ZN VDD P l=0.183881u w=2.01u 
MM20 VDD 3 ZN VDD P l=0.18516u w=2.035u 
MM19 ZN 3 VDD VDD P l=0.18u w=1.94u 
MM18 VDD B 5 VDD P l=0.18u w=0.5u 
MM17 VDD 5 2 VDD P l=0.186679u w=1.096u 
MM16 VDD 6 2 VDD P l=0.18u w=1.03u 
MM15 2 A VDD VDD P l=0.186207u w=1.102u 
MM14 VDD C2 6 VDD P l=0.18u w=1.08u 
MM13 VDD C3 6 VDD P l=0.18u w=1.15u 
MM12 VDD C1 6 VDD P l=0.18u w=1.15u 
MM11 3 2 VSS VSS N l=0.186867u w=1.066u 
MM10 VSS 3 ZN VSS N l=0.188286u w=1.383u 
MM9 ZN 3 VSS VSS N l=0.185097u w=1.342u 
MM8 ZN 3 VSS VSS N l=0.18u w=1.28u 
MM7 14 5 13 VSS N l=0.18u w=0.98u 
MM6 VSS 6 13 VSS N l=0.18u w=0.98u 
MM5 2 A 14 VSS N l=0.18u w=0.98u 
MM4 15 C2 16 VSS N l=0.18u w=0.98u 
MM3 15 C3 VSS VSS N l=0.18u w=0.98u 
MM2 6 C1 16 VSS N l=0.18u w=0.98u 
MM1 VSS B 5 VSS N l=0.18u w=0.48u 
.ENDS oaim3m11d4

.SUBCKT oan211d1 ZN  A B C1 C2 VDD VSS
MM8 ZN A 6 VDD P l=0.18u w=1.33u 
MM7 VDD B 6 VDD P l=0.184914u w=1.392u 
MM6 10 C2 VDD VDD P l=0.18u w=1.33u 
MM5 10 C1 6 VDD P l=0.18u w=1.33u 
MM4 ZN A VSS VSS N l=0.187638u w=1.084u 
MM3 8 B ZN VSS N l=0.18u w=1.01u 
MM2 8 C2 VSS VSS N l=0.186381u w=1.072u 
MM1 8 C1 VSS VSS N l=0.186502u w=1.052u 
.ENDS oan211d1

.SUBCKT oan211d2 ZN  A B C1 C2 VDD VSS
MM14 6 A 11 VDD P l=0.18u w=1.33u 
MM13 VDD B 11 VDD P l=0.184914u w=1.392u 
MM12 12 C2 VDD VDD P l=0.18u w=1.33u 
MM11 12 C1 11 VDD P l=0.18u w=1.33u 
MM10 7 6 VDD VDD P l=0.185097u w=1.342u 
MM9 ZN 7 VDD VDD P l=0.184554u w=1.502u 
MM8 VDD 7 ZN VDD P l=0.184554u w=1.502u 
MM7 6 A VSS VSS N l=0.187638u w=1.084u 
MM6 10 B 6 VSS N l=0.18u w=1.01u 
MM5 10 C2 VSS VSS N l=0.186381u w=1.072u 
MM4 10 C1 VSS VSS N l=0.186502u w=1.052u 
MM3 VSS 6 7 VSS N l=0.186381u w=1.072u 
MM2 VSS 7 ZN VSS N l=0.186826u w=1.002u 
MM1 VSS 7 ZN VSS N l=0.186826u w=1.002u 
.ENDS oan211d2

.SUBCKT oan211d4 ZN  A B C1 C2 VDD VSS
MM16 3 2 VDD VDD P l=0.185097u w=1.342u 
MM14 VDD 3 ZN VDD P l=0.183486u w=1.962u 
MM15 ZN 3 VDD VDD P l=0.183333u w=2.052u 
MM13 ZN 3 VDD VDD P l=0.18u w=1.99u 
MM12 2 A 11 VDD P l=0.18u w=1.33u 
MM11 VDD B 11 VDD P l=0.184914u w=1.392u 
MM10 12 C2 VDD VDD P l=0.18u w=1.33u 
MM9 12 C1 11 VDD P l=0.18u w=1.33u 
MM8 VSS 2 3 VSS N l=0.186381u w=1.072u 
MM7 ZN 3 VSS VSS N l=0.184465u w=1.532u 
MM5 VSS 3 ZN VSS N l=0.18u w=0.94u 
MM6 VSS 3 ZN VSS N l=0.184465u w=1.532u 
MM4 2 A VSS VSS N l=0.187638u w=1.084u 
MM3 10 B 2 VSS N l=0.18u w=1.01u 
MM2 10 C2 VSS VSS N l=0.186381u w=1.072u 
MM1 10 C1 VSS VSS N l=0.186502u w=1.052u 
.ENDS oan211d4

.SUBCKT or02d0 Z  A1 A2 VDD VSS
MM5 VDD 3 Z VDD P l=0.18u w=0.75u 
MM6 7 A2 VDD VDD P l=0.18u w=0.89u 
MM4 3 A1 7 VDD P l=0.18u w=0.89u 
MM2 Z 3 VSS VSS N l=0.18u w=0.5u 
MM3 VSS A2 3 VSS N l=0.18u w=0.48u 
MM1 VSS A1 3 VSS N l=0.18u w=0.48u 
.ENDS or02d0

.SUBCKT or02d1 Z  A1 A2 VDD VSS
MM5 Z 3 VDD VDD P l=0.18u w=1.5u 
MM6 7 A2 VDD VDD P l=0.18u w=0.89u 
MM4 3 A1 7 VDD P l=0.18u w=0.89u 
MM2 Z 3 VSS VSS N l=0.18u w=1u 
MM3 VSS A2 3 VSS N l=0.18u w=0.48u 
MM1 VSS A1 3 VSS N l=0.18u w=0.48u 
.ENDS or02d1

.SUBCKT or02d2 Z  A1 A2 VDD VSS
MM8 VDD 2 Z VDD P l=0.187239u w=1.583u 
MM7 Z 2 VDD VDD P l=0.18u w=1.48u 
MM6 7 A2 VDD VDD P l=0.18u w=0.89u 
MM5 2 A1 7 VDD P l=0.18u w=0.89u 
MM4 VSS 2 Z VSS N l=0.186502u w=1.052u 
MM3 Z 2 VSS VSS N l=0.18u w=0.99u 
MM2 VSS A2 2 VSS N l=0.18u w=0.48u 
MM1 VSS A1 2 VSS N l=0.18u w=0.48u 
.ENDS or02d2

.SUBCKT or02d4 Z  A1 A2 VDD VSS
MM9 VDD 2 Z VDD P l=0.183417u w=2.002u 
MM10 Z 2 VDD VDD P l=0.183417u w=2.002u 
MM8 Z 2 VDD VDD P l=0.183417u w=2.002u 
MM7 VDD A2 7 VDD P l=0.18u w=0.89u 
MM6 2 A1 7 VDD P l=0.18u w=0.89u 
MM5 Z 2 VSS VSS N l=0.185135u w=1.332u 
MM4 Z 2 VSS VSS N l=0.185135u w=1.332u 
MM3 Z 2 VSS VSS N l=0.185135u w=1.332u 
MM2 VSS A2 2 VSS N l=0.18u w=0.48u 
MM1 VSS A1 2 VSS N l=0.18u w=0.48u 
.ENDS or02d4

.SUBCKT or03d0 Z  A1 A2 A3 VDD VSS
MM7 Z 3 VDD VDD P l=0.18u w=1u 
MM8 8 A3 VDD VDD P l=0.18u w=1u 
MM6 8 A2 9 VDD P l=0.18u w=1u 
MM5 3 A1 9 VDD P l=0.18u w=1u 
MM3 VSS 3 Z VSS N l=0.18u w=0.67u 
MM4 VSS A3 3 VSS N l=0.18u w=0.5u 
MM2 VSS A2 3 VSS N l=0.18u w=0.5u 
MM1 VSS A1 3 VSS N l=0.18u w=0.5u 
.ENDS or03d0

.SUBCKT or03d1 Z  A1 A2 A3 VDD VSS
MM7 Z 3 VDD VDD P l=0.18u w=1.5u 
MM8 8 A3 VDD VDD P l=0.18u w=1u 
MM6 8 A2 9 VDD P l=0.18u w=1u 
MM5 3 A1 9 VDD P l=0.18u w=1u 
MM3 VSS 3 Z VSS N l=0.18u w=1u 
MM4 VSS A3 3 VSS N l=0.18u w=0.5u 
MM2 VSS A2 3 VSS N l=0.18u w=0.5u 
MM1 VSS A1 3 VSS N l=0.18u w=0.5u 
.ENDS or03d1

.SUBCKT or03d2 Z  A1 A2 A3 VDD VSS
MM10 Z 2 VDD VDD P l=0.185u w=1.502u 
MM9 Z 2 VDD VDD P l=0.185u w=1.506u 
MM8 8 A3 VDD VDD P l=0.18u w=1u 
MM7 8 A2 9 VDD P l=0.18u w=1u 
MM6 2 A1 9 VDD P l=0.18u w=1u 
MM5 VSS 2 Z VSS N l=0.187u w=1.006u 
MM4 Z 2 VSS VSS N l=0.187u w=1.002u 
MM3 VSS A3 2 VSS N l=0.18u w=0.5u 
MM2 VSS A2 2 VSS N l=0.18u w=0.5u 
MM1 VSS A1 2 VSS N l=0.18u w=0.5u 
.ENDS or03d2

.SUBCKT or03d4 Z  A1 A2 A3 VDD VSS
MM12 Z 2 VDD VDD P l=0.183881u w=2.01u 
MM11 Z 2 VDD VDD P l=0.18516u w=2.035u 
MM10 Z 2 VDD VDD P l=0.18u w=1.94u 
MM9 8 A3 VDD VDD P l=0.18u w=0.98u 
MM8 8 A2 9 VDD P l=0.18u w=0.98u 
MM7 2 A1 9 VDD P l=0.18u w=0.98u 
MM5 VSS 2 Z VSS N l=0.185778u w=1.35u 
MM6 VSS 2 Z VSS N l=0.186451u w=1.358u 
MM4 VSS 2 Z VSS N l=0.18u w=1.28u 
MM3 VSS A3 2 VSS N l=0.18u w=0.49u 
MM2 2 A2 VSS VSS N l=0.18u w=0.49u 
MM1 2 A1 VSS VSS N l=0.18u w=0.49u 
.ENDS or03d4

.SUBCKT or04d0 Z  A1 A2 A3 A4 VDD VSS
MM10 VDD 2 Z VDD P l=0.18u w=0.75u 
MM9 VDD A4 9 VDD P l=0.18527u w=1.48u 
MM8 10 A3 9 VDD P l=0.18u w=1.41u 
MM7 10 A2 11 VDD P l=0.18u w=1.41u 
MM6 2 A1 11 VDD P l=0.18u w=1.41u 
MM5 VSS 2 Z VSS N l=0.18u w=0.5u 
MM4 VSS A4 2 VSS N l=0.18u w=0.62u 
MM3 VSS A3 2 VSS N l=0.18u w=0.62u 
MM2 VSS A2 2 VSS N l=0.18u w=0.48u 
MM1 VSS A1 2 VSS N l=0.18u w=0.48u 
.ENDS or04d0

.SUBCKT or04d1 Z  A1 A2 A3 A4 VDD VSS
MM9 VDD 3 Z VDD P l=0.18u w=1.5u 
MM10 VDD A4 9 VDD P l=0.18527u w=1.48u 
MM8 10 A3 9 VDD P l=0.18u w=1.41u 
MM7 11 A2 10 VDD P l=0.18u w=1.41u 
MM6 11 A1 3 VDD P l=0.18u w=1.41u 
MM4 Z 3 VSS VSS N l=0.18u w=1u 
MM5 VSS A4 3 VSS N l=0.18u w=0.62u 
MM3 VSS A3 3 VSS N l=0.18u w=0.62u 
MM2 VSS A2 3 VSS N l=0.18u w=0.48u 
MM1 VSS A1 3 VSS N l=0.18u w=0.48u 
.ENDS or04d1

.SUBCKT or04d2 Z  A1 A2 A3 A4 VDD VSS
MM11 VDD 3 Z VDD P l=0.184554u w=1.502u 
MM10 VDD 3 Z VDD P l=0.184554u w=1.502u 
MM12 VDD A4 9 VDD P l=0.18527u w=1.48u 
MM9 10 A3 9 VDD P l=0.18u w=1.41u 
MM8 11 A2 10 VDD P l=0.18u w=1.41u 
MM7 11 A1 3 VDD P l=0.18u w=1.41u 
MM5 Z 3 VSS VSS N l=0.186826u w=1.002u 
MM4 Z 3 VSS VSS N l=0.186826u w=1.002u 
MM6 VSS A4 3 VSS N l=0.18u w=0.62u 
MM3 VSS A3 3 VSS N l=0.18u w=0.62u 
MM2 VSS A2 3 VSS N l=0.18u w=0.48u 
MM1 VSS A1 3 VSS N l=0.18u w=0.48u 
.ENDS or04d2

.SUBCKT or04d4 Z  A1 A2 A3 A4 VDD VSS
MM12 Z 3 VDD VDD P l=0.183417u w=2.002u 
MM13 VDD 3 Z VDD P l=0.183417u w=2.002u 
MM11 VDD 3 Z VDD P l=0.183417u w=2.002u 
MM14 VDD A4 9 VDD P l=0.18527u w=1.48u 
MM10 10 A3 9 VDD P l=0.18u w=1.41u 
MM9 11 A2 10 VDD P l=0.18u w=1.41u 
MM8 11 A1 3 VDD P l=0.18u w=1.41u 
MM6 Z 3 VSS VSS N l=0.185135u w=1.332u 
MM5 Z 3 VSS VSS N l=0.185135u w=1.332u 
MM4 Z 3 VSS VSS N l=0.185135u w=1.332u 
MM7 VSS A4 3 VSS N l=0.18u w=0.62u 
MM3 VSS A3 3 VSS N l=0.18u w=0.62u 
MM2 VSS A2 3 VSS N l=0.18u w=0.48u 
MM1 VSS A1 3 VSS N l=0.18u w=0.48u 
.ENDS or04d4

.SUBCKT ora211d1 Z  A B C1 C2 VDD VSS
MM9 VDD 3 Z VDD P l=0.1852u w=1.5u 
MM8 3 A VDD VDD P l=0.18u w=0.81u 
MM7 VDD B 3 VDD P l=0.18u w=0.82u 
MM6 11 C1 3 VDD P l=0.18u w=1.45u 
MM10 11 C2 VDD VDD P l=0.18u w=1.45u 
MM5 8 C2 VSS VSS N l=0.18u w=0.75u 
MM4 Z 3 VSS VSS N l=0.18u w=1u 
MM3 3 A 10 VSS N l=0.18u w=0.99u 
MM2 8 B 10 VSS N l=0.18u w=0.99u 
MM1 VSS C1 8 VSS N l=0.187358u w=1.06u 
.ENDS ora211d1

.SUBCKT ora211d2 Z  A B C1 C2 VDD VSS
MM11 VDD 3 Z VDD P l=0.18u w=1.5u 
MM10 Z 3 VDD VDD P l=0.18u w=1.5u 
MM9 VDD B 3 VDD P l=0.18u w=0.82u 
MM7 11 C1 3 VDD P l=0.18u w=1.45u 
MM8 VDD A 3 VDD P l=0.18u w=0.82u 
MM12 11 C2 VDD VDD P l=0.18u w=1.45u 
MM6 VSS C2 9 VSS N l=0.18u w=0.75u 
MM5 Z 3 VSS VSS N l=0.186998u w=1.046u 
MM4 Z 3 VSS VSS N l=0.18u w=0.98u 
MM3 9 B 10 VSS N l=0.18u w=0.99u 
MM2 3 A 10 VSS N l=0.18u w=0.99u 
MM1 VSS C1 9 VSS N l=0.187358u w=1.06u 
.ENDS ora211d2

.SUBCKT ora211d4 Z  A B C1 C2 VDD VSS
MM14 VDD C2 11 VDD P l=0.18u w=1.45u 
MM8 3 C1 11 VDD P l=0.18u w=1.45u 
MM13 Z 3 VDD VDD P l=0.183861u w=2.02u 
MM12 Z 3 VDD VDD P l=0.185134u w=2.045u 
MM11 VDD 3 Z VDD P l=0.18u w=1.95u 
MM10 VDD A 3 VDD P l=0.18u w=0.81u 
MM9 VDD B 3 VDD P l=0.18u w=0.82u 
MM7 VSS C2 8 VSS N l=0.18u w=0.75u 
MM6 Z 3 VSS VSS N l=0.188286u w=1.383u 
MM5 VSS 3 Z VSS N l=0.185438u w=1.346u 
MM4 Z 3 VSS VSS N l=0.18u w=1.28u 
MM3 3 A 10 VSS N l=0.18u w=0.99u 
MM2 8 B 10 VSS N l=0.18u w=0.99u 
MM1 8 C1 VSS VSS N l=0.18u w=1.07u 
.ENDS ora211d4

.SUBCKT ora21d1 Z  A B1 B2 VDD VSS
MM7 VDD 3 Z VDD P l=0.18u w=1.5u 
MM6 VDD A 3 VDD P l=0.18u w=0.9u 
MM5 3 B1 9 VDD P l=0.18u w=1.51u 
MM8 VDD B2 9 VDD P l=0.18u w=1.51u 
MM4 7 B2 VSS VSS N l=0.186142u w=1.27u 
MM3 7 A 3 VSS N l=0.185787u w=1.182u 
MM2 7 B1 VSS VSS N l=0.185787u w=1.182u 
MM1 Z 3 VSS VSS N l=0.1878u w=1u 
.ENDS ora21d1

.SUBCKT ora21d2 Z  A B1 B2 VDD VSS
MM10 Z 2 VDD VDD P l=0.184465u w=1.532u 
MM9 Z 2 VDD VDD P l=0.18u w=1.47u 
MM8 VDD A 2 VDD P l=0.18u w=0.9u 
MM6 2 B1 9 VDD P l=0.18u w=1.51u 
MM7 VDD B2 9 VDD P l=0.18u w=1.51u 
MM5 7 A 2 VSS N l=0.185787u w=1.182u 
MM4 7 B2 VSS VSS N l=0.186142u w=1.27u 
MM3 7 B1 VSS VSS N l=0.185787u w=1.182u 
MM2 Z 2 VSS VSS N l=0.1878u w=1u 
MM1 Z 2 VSS VSS N l=0.1878u w=1u 
.ENDS ora21d2

.SUBCKT ora21d4 Z  A B1 B2 VDD VSS
MM11 Z 2 VDD VDD P l=0.183417u w=2.002u 
MM12 VDD 2 Z VDD P l=0.183417u w=2.002u 
MM10 VDD 2 Z VDD P l=0.183417u w=2.002u 
MM9 VDD A 2 VDD P l=0.18u w=0.9u 
MM7 2 B1 9 VDD P l=0.18u w=1.51u 
MM8 VDD B2 9 VDD P l=0.18u w=1.51u 
MM6 Z 2 VSS VSS N l=0.185135u w=1.332u 
MM5 Z 2 VSS VSS N l=0.185135u w=1.332u 
MM4 Z 2 VSS VSS N l=0.185135u w=1.332u 
MM3 8 A 2 VSS N l=0.185787u w=1.182u 
MM2 8 B2 VSS VSS N l=0.186142u w=1.27u 
MM1 8 B1 VSS VSS N l=0.185787u w=1.182u 
.ENDS ora21d4

.SUBCKT ora311d1 Z  A B C1 C2 C3 VDD VSS
MM11 Z 3 VDD VDD P l=0.18u w=1.5u 
MM12 12 C2 13 VDD P l=0.18u w=1.5u 
MM10 12 C3 VDD VDD P l=0.18u w=1.5u 
MM9 3 A VDD VDD P l=0.186867u w=1.066u 
MM8 13 C1 3 VDD P l=0.18u w=1.5u 
MM7 VDD B 3 VDD P l=0.186693u w=1.022u 
MM5 Z 3 VSS VSS N l=0.18u w=1u 
MM6 VSS C2 9 VSS N l=0.186207u w=1.102u 
MM4 VSS C3 9 VSS N l=0.18u w=1.04u 
MM3 11 A 3 VSS N l=0.18u w=0.79u 
MM2 VSS C1 9 VSS N l=0.186693u w=1.022u 
MM1 9 B 11 VSS N l=0.18u w=0.79u 
.ENDS ora311d1

.SUBCKT ora311d2 Z  A B C1 C2 C3 VDD VSS
MM14 Z 2 VDD VDD P l=0.184554u w=1.502u 
MM13 VDD 2 Z VDD P l=0.184861u w=1.506u 
MM11 2 A VDD VDD P l=0.186803u w=1.076u 
MM12 12 C3 VDD VDD P l=0.18u w=1.49u 
MM10 12 C2 13 VDD P l=0.18u w=1.49u 
MM9 13 C1 2 VDD P l=0.18u w=1.49u 
MM8 VDD B 2 VDD P l=0.186759u w=1.012u 
MM7 Z 2 VSS VSS N l=0.187276u w=1.006u 
MM6 VSS 2 Z VSS N l=0.186826u w=1.002u 
MM4 11 A 2 VSS N l=0.18u w=0.79u 
MM5 VSS C3 9 VSS N l=0.18u w=1.04u 
MM3 VSS C2 9 VSS N l=0.186207u w=1.102u 
MM2 VSS C1 9 VSS N l=0.186693u w=1.022u 
MM1 9 B 11 VSS N l=0.18u w=0.79u 
.ENDS ora311d2

.SUBCKT ora311d4 Z  A B C1 C2 C3 VDD VSS
MM15 Z 3 VDD VDD P l=0.183881u w=2.01u 
MM14 Z 3 VDD VDD P l=0.18516u w=2.035u 
MM13 VDD 3 Z VDD P l=0.18u w=1.94u 
MM12 3 A VDD VDD P l=0.186867u w=1.066u 
MM16 12 C3 VDD VDD P l=0.18u w=1.49u 
MM11 12 C2 13 VDD P l=0.18u w=1.49u 
MM10 13 C1 3 VDD P l=0.18u w=1.49u 
MM9 VDD B 3 VDD P l=0.18u w=0.95u 
MM7 Z 3 VSS VSS N l=0.188286u w=1.383u 
MM6 VSS 3 Z VSS N l=0.185097u w=1.342u 
MM5 Z 3 VSS VSS N l=0.18u w=1.28u 
MM4 11 A 3 VSS N l=0.18u w=0.79u 
MM8 VSS C3 10 VSS N l=0.18u w=1.04u 
MM3 VSS C2 10 VSS N l=0.186207u w=1.102u 
MM2 VSS C1 10 VSS N l=0.186693u w=1.022u 
MM1 10 B 11 VSS N l=0.18u w=0.79u 
.ENDS ora311d4

.SUBCKT ora31d1 Z  A B1 B2 B3 VDD VSS
MM9 VDD 3 Z VDD P l=0.18u w=1.5u 
MM10 11 B2 10 VDD P l=0.18u w=1.62u 
MM8 VDD B3 10 VDD P l=0.18u w=1.62u 
MM7 VDD A 3 VDD P l=0.188235u w=1.122u 
MM6 11 B1 3 VDD P l=0.18u w=1.62u 
MM5 VSS B2 8 VSS N l=0.18u w=1.07u 
MM3 VSS B3 8 VSS N l=0.18u w=1.07u 
MM4 Z 3 VSS VSS N l=0.186826u w=1.002u 
MM2 8 A 3 VSS N l=0.18u w=0.9u 
MM1 VSS B1 8 VSS N l=0.186501u w=1.126u 
.ENDS ora31d1

.SUBCKT ora31d2 Z  A B1 B2 B3 VDD VSS
MM12 VDD 2 Z VDD P l=0.185662u w=1.632u 
MM11 VDD 2 Z VDD P l=0.18u w=1.55u 
MM10 VDD B3 10 VDD P l=0.18u w=1.62u 
MM8 11 B2 10 VDD P l=0.18u w=1.62u 
MM9 VDD A 2 VDD P l=0.188235u w=1.122u 
MM7 11 B1 2 VDD P l=0.18u w=1.62u 
MM6 Z 2 VSS VSS N l=0.187358u w=1.06u 
MM5 Z 2 VSS VSS N l=0.186502u w=1.052u 
MM4 8 B3 VSS VSS N l=0.18u w=1.07u 
MM2 VSS B2 8 VSS N l=0.18u w=1.07u 
MM3 8 A 2 VSS N l=0.18u w=0.9u 
MM1 VSS B1 8 VSS N l=0.186501u w=1.126u 
.ENDS ora31d2

.SUBCKT ora31d4 Z  A B1 B2 B3 VDD VSS
MM12 VDD 3 Z VDD P l=0.184845u w=1.808u 
MM11 VDD 3 Z VDD P l=0.18u w=1.73u 
MM10 VDD 3 Z VDD P l=0.18459u w=1.804u 
MM13 VDD B3 10 VDD P l=0.18u w=1.62u 
MM8 11 B2 10 VDD P l=0.18u w=1.62u 
MM9 VDD A 3 VDD P l=0.188235u w=1.122u 
MM7 11 B1 3 VDD P l=0.18u w=1.62u 
MM6 VSS B3 9 VSS N l=0.18u w=1.07u 
MM2 VSS B2 9 VSS N l=0.18u w=1.07u 
MM5 Z 3 VSS VSS N l=0.190556u w=1.779u 
MM4 Z 3 VSS VSS N l=0.19031u w=1.775u 
MM3 9 A 3 VSS N l=0.18u w=0.9u 
MM1 VSS B1 9 VSS N l=0.186501u w=1.126u 
.ENDS ora31d4

.SUBCKT sdbrb1 Q QN  CDN CP D SC SD SDN VDD VSS
MM43 11 SC VDD VDD P l=0.18u w=0.95u 
MM42 VDD 7 8 VDD P l=0.18u w=0.52u 
MM41 23 8 VDD VDD P l=0.18u w=0.52u 
MM38 23 11 24 VDD P l=0.18u w=0.52u 
MM40 25 9 24 VDD P l=0.18u w=0.52u 
MM39 VDD D 25 VDD P l=0.18u w=0.52u 
MM37 VDD 11 9 VDD P l=0.18u w=0.5u 
MM26 3 CP VDD VDD P l=0.18u w=0.97u 
MM25 VDD SD 7 VDD P l=0.18u w=0.52u 
MM48 IPM 2 24 VDD P l=0.18u w=0.6u 
MM47 IPM 3 18 VDD P l=0.18u w=0.6u 
MM34 15 IPM VDD VDD P l=0.18u w=0.86u 
MM35 22 2 IPS VDD P l=0.18u w=0.76u 
MM32 22 SDN VDD VDD P l=0.186264u w=1.092u 
MM31 VDD SDN 15 VDD P l=0.186502u w=1.052u 
MM30 IPS 3 15 VDD P l=0.18u w=0.76u 
MM29 18 15 VDD VDD P l=0.18u w=0.6u 
MM28 18 CDN VDD VDD P l=0.18u w=0.6u 
MM27 2 3 VDD VDD P l=0.18u w=0.76u 
MM45 QN IPS VDD VDD P l=0.18u w=1.5u 
MM46 VDD IPS 12 VDD P l=0.186115u w=1.354u 
MM44 12 CDN VDD VDD P l=0.18u w=1.28u 
MM36 VDD 12 Q VDD P l=0.18u w=1.5u 
MM33 22 12 VDD VDD P l=0.186264u w=1.092u 
MM24 18 2 IPM VSS N l=0.18u w=0.44u 
MM22 IPM 3 24 VSS N l=0.18u w=0.44u 
MM23 15 2 IPS VSS N l=0.18u w=0.6u 
MM21 22 3 IPS VSS N l=0.18u w=0.6u 
MM17 26 SDN 22 VSS N l=0.18u w=0.8u 
MM19 VSS 12 26 VSS N l=0.18u w=0.8u 
MM16 27 SDN 15 VSS N l=0.18u w=0.75u 
MM20 27 IPM VSS VSS N l=0.18u w=0.75u 
MM14 18 CDN 28 VSS N l=0.18u w=0.75u 
MM15 28 15 VSS VSS N l=0.18u w=0.75u 
MM13 29 CDN 12 VSS N l=0.18u w=1.21u 
MM18 VSS IPS 29 VSS N l=0.18u w=1.21u 
MM12 Q 12 VSS VSS N l=0.18u w=1.08u 
MM11 QN IPS VSS VSS N l=0.18u w=1.08u 
MM10 8 7 VSS VSS N l=0.18u w=0.48u 
MM9 23 8 VSS VSS N l=0.18u w=0.48u 
MM8 23 9 24 VSS N l=0.18u w=0.48u 
MM6 VSS 11 9 VSS N l=0.18u w=0.43u 
MM5 24 11 25 VSS N l=0.18u w=0.48u 
MM7 VSS D 25 VSS N l=0.18u w=0.48u 
MM2 VSS SD 7 VSS N l=0.18u w=0.43u 
MM4 2 3 VSS VSS N l=0.18u w=0.52u 
MM3 VSS CP 3 VSS N l=0.18u w=0.52u 
MM1 11 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdbrb1

.SUBCKT sdbrb2 Q QN  CDN CP D SC SD SDN VDD VSS
MM33 22 6 VDD VDD P l=0.186264u w=1.092u 
MM29 2 3 VDD VDD P l=0.18u w=0.76u 
MM42 13 SC VDD VDD P l=0.18u w=0.95u 
MM41 VDD 9 10 VDD P l=0.18u w=0.52u 
MM40 23 10 VDD VDD P l=0.18u w=0.52u 
MM37 23 13 24 VDD P l=0.18u w=0.52u 
MM39 25 11 24 VDD P l=0.18u w=0.52u 
MM38 VDD D 25 VDD P l=0.18u w=0.52u 
MM36 VDD 13 11 VDD P l=0.18u w=0.5u 
MM28 3 CP VDD VDD P l=0.18u w=0.97u 
MM27 VDD SD 9 VDD P l=0.18u w=0.52u 
MM52 IPM 2 24 VDD P l=0.18u w=0.6u 
MM51 IPM 3 18 VDD P l=0.18u w=0.6u 
MM50 18 4 VDD VDD P l=0.18u w=0.6u 
MM49 18 CDN VDD VDD P l=0.18u w=0.6u 
MM34 VDD IPM 4 VDD P l=0.18u w=0.86u 
MM35 22 2 IPS VDD P l=0.18u w=0.76u 
MM32 22 SDN VDD VDD P l=0.186264u w=1.092u 
MM31 VDD SDN 4 VDD P l=0.186502u w=1.052u 
MM30 IPS 3 4 VDD P l=0.18u w=0.76u 
MM48 VDD 6 Q VDD P l=0.184845u w=1.61u 
MM47 VDD 6 Q VDD P l=0.18u w=1.54u 
MM45 QN IPS VDD VDD P l=0.18u w=1.54u 
MM44 VDD IPS QN VDD P l=0.18513u w=1.614u 
MM46 VDD IPS 6 VDD P l=0.186115u w=1.354u 
MM43 6 CDN VDD VDD P l=0.18u w=1.28u 
MM26 18 2 IPM VSS N l=0.18u w=0.44u 
MM24 IPM 3 24 VSS N l=0.18u w=0.44u 
MM25 4 2 IPS VSS N l=0.18u w=0.6u 
MM23 22 3 IPS VSS N l=0.18u w=0.6u 
MM19 26 SDN 22 VSS N l=0.18u w=0.8u 
MM21 VSS 6 26 VSS N l=0.18u w=0.8u 
MM18 27 SDN 4 VSS N l=0.18u w=0.75u 
MM22 27 IPM VSS VSS N l=0.18u w=0.75u 
MM16 18 CDN 28 VSS N l=0.18u w=0.75u 
MM17 28 4 VSS VSS N l=0.18u w=0.75u 
MM15 29 CDN 6 VSS N l=0.18u w=1.21u 
MM20 VSS IPS 29 VSS N l=0.18u w=1.21u 
MM14 10 9 VSS VSS N l=0.18u w=0.48u 
MM13 23 10 VSS VSS N l=0.18u w=0.48u 
MM12 23 11 24 VSS N l=0.18u w=0.48u 
MM10 VSS 13 11 VSS N l=0.18u w=0.43u 
MM9 24 13 25 VSS N l=0.18u w=0.48u 
MM11 VSS D 25 VSS N l=0.18u w=0.48u 
MM6 VSS SD 9 VSS N l=0.18u w=0.43u 
MM8 2 3 VSS VSS N l=0.18u w=0.52u 
MM7 VSS CP 3 VSS N l=0.18u w=0.52u 
MM5 Q 6 VSS VSS N l=0.186502u w=1.052u 
MM4 Q 6 VSS VSS N l=0.186502u w=1.052u 
MM3 VSS IPS QN VSS N l=0.186502u w=1.052u 
MM2 QN IPS VSS VSS N l=0.186502u w=1.052u 
MM1 13 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdbrb2

.SUBCKT sdcfq1 Q  CDN CPN D SC SD VDD VSS
MM41 VDD 3 19 VDD P l=0.18u w=0.55u 
MM35 19 CDN VDD VDD P l=0.18u w=0.52u 
MM42 21 2 IPS VDD P l=0.18u w=0.75u 
MM40 VDD 4 21 VDD P l=0.18u w=0.71u 
MM37 VDD 4 Q VDD P l=0.184524u w=1.512u 
MM38 4 IPS VDD VDD P l=0.185479u w=1.336u 
MM36 VDD CDN 4 VDD P l=0.18u w=1.27u 
MM34 IPS 8 3 VDD P l=0.18u w=0.75u 
MM39 VDD IPM 3 VDD P l=0.18u w=0.75u 
MM33 VDD 9 10 VDD P l=0.18u w=0.52u 
MM32 22 10 VDD VDD P l=0.18u w=0.52u 
MM29 22 13 17 VDD P l=0.18u w=0.58u 
MM31 23 11 17 VDD P l=0.18u w=0.42u 
MM30 VDD D 23 VDD P l=0.18u w=0.52u 
MM28 VDD 13 11 VDD P l=0.18u w=0.52u 
MM27 IPM 2 17 VDD P l=0.18u w=0.6u 
MM26 IPM 8 19 VDD P l=0.18u w=0.6u 
MM25 8 2 VDD VDD P l=0.18u w=0.68u 
MM24 2 CPN VDD VDD P l=0.18u w=0.68u 
MM23 VDD SD 9 VDD P l=0.18u w=0.52u 
MM22 13 SC VDD VDD P l=0.18u w=0.52u 
MM21 17 8 IPM VSS N l=0.18u w=0.44u 
MM19 IPM 2 19 VSS N l=0.18u w=0.44u 
MM18 3 2 IPS VSS N l=0.18u w=0.6u 
MM15 3 IPM VSS VSS N l=0.18u w=0.52u 
MM20 21 8 IPS VSS N l=0.18u w=0.6u 
MM16 21 4 VSS VSS N l=0.18u w=0.6u 
MM13 24 CDN 19 VSS N l=0.18u w=0.75u 
MM17 VSS 3 24 VSS N l=0.18u w=0.75u 
MM12 4 CDN 25 VSS N l=0.18u w=1.11u 
MM14 VSS IPS 25 VSS N l=0.18u w=1.11u 
MM11 10 9 VSS VSS N l=0.18u w=0.42u 
MM10 22 10 VSS VSS N l=0.18u w=0.44u 
MM9 22 11 17 VSS N l=0.18u w=0.44u 
MM7 VSS 13 11 VSS N l=0.18u w=0.43u 
MM6 17 13 23 VSS N l=0.18u w=0.44u 
MM8 VSS D 23 VSS N l=0.18u w=0.44u 
MM3 VSS SD 9 VSS N l=0.18u w=0.43u 
MM5 8 2 VSS VSS N l=0.18u w=0.52u 
MM4 VSS CPN 2 VSS N l=0.18u w=0.52u 
MM2 VSS 4 Q VSS N l=0.186441u w=1.062u 
MM1 13 SC VSS VSS N l=0.18u w=0.43u 
.ENDS sdcfq1

.SUBCKT sdcfq2 Q  CDN CPN D SC SD VDD VSS
MM43 IPM 2 17 VDD P l=0.18u w=0.6u 
MM42 IPM 3 19 VDD P l=0.18u w=0.6u 
MM40 VDD 4 19 VDD P l=0.18u w=0.55u 
MM33 19 CDN VDD VDD P l=0.18u w=0.52u 
MM41 21 2 IPS VDD P l=0.18u w=0.75u 
MM39 VDD 5 21 VDD P l=0.18u w=0.71u 
MM36 VDD 5 Q VDD P l=0.184494u w=1.522u 
MM35 Q 5 VDD VDD P l=0.184494u w=1.522u 
MM37 VDD IPS 5 VDD P l=0.184797u w=1.526u 
MM34 VDD CDN 5 VDD P l=0.18u w=1.46u 
MM32 IPS 3 4 VDD P l=0.18u w=0.75u 
MM38 VDD IPM 4 VDD P l=0.18u w=0.75u 
MM31 VDD 9 10 VDD P l=0.18u w=0.52u 
MM30 22 10 VDD VDD P l=0.18u w=0.52u 
MM27 22 13 17 VDD P l=0.18u w=0.58u 
MM29 23 11 17 VDD P l=0.18u w=0.42u 
MM28 VDD D 23 VDD P l=0.18u w=0.52u 
MM26 VDD 13 11 VDD P l=0.18u w=0.52u 
MM25 3 2 VDD VDD P l=0.18u w=0.68u 
MM24 2 CPN VDD VDD P l=0.18u w=0.68u 
MM23 VDD SD 9 VDD P l=0.18u w=0.52u 
MM22 13 SC VDD VDD P l=0.18u w=0.52u 
MM21 17 3 IPM VSS N l=0.18u w=0.44u 
MM19 IPM 2 19 VSS N l=0.18u w=0.44u 
MM18 4 2 IPS VSS N l=0.18u w=0.6u 
MM15 4 IPM VSS VSS N l=0.18u w=0.52u 
MM20 21 3 IPS VSS N l=0.18u w=0.6u 
MM16 21 5 VSS VSS N l=0.18u w=0.6u 
MM13 5 CDN 24 VSS N l=0.18u w=1.3u 
MM14 VSS IPS 24 VSS N l=0.18u w=1.3u 
MM12 25 CDN 19 VSS N l=0.18u w=0.75u 
MM17 VSS 4 25 VSS N l=0.18u w=0.75u 
MM11 VSS 5 Q VSS N l=0.184132u w=2.004u 
MM10 10 9 VSS VSS N l=0.18u w=0.42u 
MM9 22 10 VSS VSS N l=0.18u w=0.44u 
MM8 22 11 17 VSS N l=0.18u w=0.44u 
MM6 VSS 13 11 VSS N l=0.18u w=0.43u 
MM5 17 13 23 VSS N l=0.18u w=0.44u 
MM7 VSS D 23 VSS N l=0.18u w=0.44u 
MM2 VSS SD 9 VSS N l=0.18u w=0.43u 
MM4 3 2 VSS VSS N l=0.18u w=0.52u 
MM3 VSS CPN 2 VSS N l=0.18u w=0.52u 
MM1 13 SC VSS VSS N l=0.18u w=0.43u 
.ENDS sdcfq2

.SUBCKT sdcrb1 Q QN  CDN CP D SC SD VDD VSS
MM44 IPM 2 23 VDD P l=0.18u w=0.6u 
MM43 IPM 3 20 VDD P l=0.18u w=0.6u 
MM41 VDD 4 20 VDD P l=0.18u w=0.55u 
MM36 20 CDN VDD VDD P l=0.18u w=0.52u 
MM42 21 2 IPS VDD P l=0.18u w=0.75u 
MM40 VDD 5 21 VDD P l=0.18u w=0.75u 
MM39 4 IPM VDD VDD P l=0.18u w=1u 
MM35 4 3 IPS VDD P l=0.18u w=0.75u 
MM38 VDD IPS 5 VDD P l=0.185875u w=1.246u 
MM37 VDD CDN 5 VDD P l=0.18u w=1.18u 
MM34 VDD 9 10 VDD P l=0.18u w=0.52u 
MM33 22 10 VDD VDD P l=0.18u w=0.52u 
MM30 22 13 23 VDD P l=0.18u w=0.52u 
MM32 24 11 23 VDD P l=0.18u w=0.52u 
MM31 VDD D 24 VDD P l=0.18u w=0.52u 
MM29 VDD 13 11 VDD P l=0.18u w=0.5u 
MM28 VDD 5 Q VDD P l=0.185342u w=1.46u 
MM27 VDD IPS QN VDD P l=0.184711u w=1.452u 
MM26 2 3 VDD VDD P l=0.18u w=0.76u 
MM25 3 CP VDD VDD P l=0.18u w=0.97u 
MM24 VDD SD 9 VDD P l=0.18u w=0.52u 
MM23 13 SC VDD VDD P l=0.18u w=0.52u 
MM22 IPM 2 20 VSS N l=0.18u w=0.44u 
MM20 23 3 IPM VSS N l=0.18u w=0.44u 
MM21 4 2 IPS VSS N l=0.18u w=0.6u 
MM19 21 3 IPS VSS N l=0.18u w=0.6u 
MM17 21 5 VSS VSS N l=0.18u w=0.6u 
MM16 4 IPM VSS VSS N l=0.18u w=0.75u 
MM14 25 CDN 20 VSS N l=0.18u w=0.75u 
MM18 VSS 4 25 VSS N l=0.18u w=0.75u 
MM13 5 CDN 26 VSS N l=0.18u w=1.21u 
MM15 VSS IPS 26 VSS N l=0.18u w=1.21u 
MM12 10 9 VSS VSS N l=0.18u w=0.48u 
MM11 22 10 VSS VSS N l=0.18u w=0.48u 
MM10 22 11 23 VSS N l=0.18u w=0.48u 
MM8 VSS 13 11 VSS N l=0.18u w=0.43u 
MM7 23 13 24 VSS N l=0.18u w=0.48u 
MM9 VSS D 24 VSS N l=0.18u w=0.48u 
MM4 VSS SD 9 VSS N l=0.18u w=0.43u 
MM6 2 3 VSS VSS N l=0.18u w=0.52u 
MM5 VSS CP 3 VSS N l=0.18u w=0.52u 
MM3 Q 5 VSS VSS N l=0.185377u w=1.272u 
MM2 QN IPS VSS VSS N l=0.185737u w=1.276u 
MM1 13 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdcrb1

.SUBCKT sdcrb2 Q QN  CDN CP D SC SD VDD VSS
MM48 IPM 2 23 VDD P l=0.18u w=0.6u 
MM47 IPM 3 20 VDD P l=0.18u w=0.6u 
MM45 VDD 4 20 VDD P l=0.18u w=0.55u 
MM36 20 CDN VDD VDD P l=0.18u w=0.52u 
MM46 21 2 IPS VDD P l=0.18u w=0.75u 
MM44 VDD 5 21 VDD P l=0.18u w=0.75u 
MM43 4 IPM VDD VDD P l=0.18u w=1u 
MM35 4 3 IPS VDD P l=0.18u w=0.75u 
MM42 VDD 5 Q VDD P l=0.18427u w=1.602u 
MM41 VDD 5 Q VDD P l=0.18427u w=1.602u 
MM40 VDD IPS QN VDD P l=0.18427u w=1.602u 
MM39 QN IPS VDD VDD P l=0.18427u w=1.602u 
MM38 VDD IPS 5 VDD P l=0.185438u w=1.346u 
MM37 VDD CDN 5 VDD P l=0.18u w=1.28u 
MM34 VDD 9 10 VDD P l=0.18u w=0.52u 
MM33 22 10 VDD VDD P l=0.18u w=0.52u 
MM30 22 13 23 VDD P l=0.18u w=0.52u 
MM32 24 11 23 VDD P l=0.18u w=0.52u 
MM31 VDD D 24 VDD P l=0.18u w=0.52u 
MM29 VDD 13 11 VDD P l=0.18u w=0.5u 
MM28 2 3 VDD VDD P l=0.18u w=0.76u 
MM27 3 CP VDD VDD P l=0.18u w=0.97u 
MM26 VDD SD 9 VDD P l=0.18u w=0.52u 
MM25 13 SC VDD VDD P l=0.18u w=0.52u 
MM24 IPM 2 20 VSS N l=0.18u w=0.44u 
MM22 23 3 IPM VSS N l=0.18u w=0.44u 
MM23 4 2 IPS VSS N l=0.18u w=0.6u 
MM21 21 3 IPS VSS N l=0.18u w=0.6u 
MM19 21 5 VSS VSS N l=0.18u w=0.6u 
MM18 4 IPM VSS VSS N l=0.18u w=0.75u 
MM16 25 CDN 20 VSS N l=0.18u w=0.75u 
MM20 VSS 4 25 VSS N l=0.18u w=0.75u 
MM15 5 CDN 26 VSS N l=0.18u w=1.21u 
MM17 VSS IPS 26 VSS N l=0.18u w=1.21u 
MM14 10 9 VSS VSS N l=0.18u w=0.48u 
MM13 22 10 VSS VSS N l=0.18u w=0.48u 
MM12 22 11 23 VSS N l=0.18u w=0.48u 
MM10 VSS 13 11 VSS N l=0.18u w=0.43u 
MM9 23 13 24 VSS N l=0.18u w=0.48u 
MM11 VSS D 24 VSS N l=0.18u w=0.48u 
MM6 VSS SD 9 VSS N l=0.18u w=0.43u 
MM8 2 3 VSS VSS N l=0.18u w=0.52u 
MM7 VSS CP 3 VSS N l=0.18u w=0.52u 
MM5 Q 5 VSS VSS N l=0.186502u w=1.052u 
MM4 Q 5 VSS VSS N l=0.186502u w=1.052u 
MM3 VSS IPS QN VSS N l=0.186502u w=1.052u 
MM2 VSS IPS QN VSS N l=0.186502u w=1.052u 
MM1 13 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdcrb2

.SUBCKT sdcrn1 QN  CDN CP D SC SD VDD VSS
MM42 VDD 2 19 VDD P l=0.18u w=0.55u 
MM36 19 CDN VDD VDD P l=0.18u w=0.52u 
MM41 VDD 3 21 VDD P l=0.18u w=0.76u 
MM40 IPS 4 21 VDD P l=0.18u w=0.88u 
MM37 VDD IPS QN VDD P l=0.184379u w=1.562u 
MM38 VDD IPS 3 VDD P l=0.186387u w=1.146u 
MM35 VDD CDN 3 VDD P l=0.18u w=1.08u 
MM34 2 8 IPS VDD P l=0.18u w=0.88u 
MM39 2 IPM VDD VDD P l=0.18u w=0.88u 
MM33 VDD 9 10 VDD P l=0.18u w=0.52u 
MM32 22 10 VDD VDD P l=0.18u w=0.52u 
MM29 22 13 17 VDD P l=0.18u w=0.52u 
MM31 23 11 17 VDD P l=0.18u w=0.52u 
MM30 VDD D 23 VDD P l=0.18u w=0.52u 
MM28 VDD 13 11 VDD P l=0.18u w=0.5u 
MM27 IPM 8 19 VDD P l=0.18u w=0.6u 
MM26 IPM 4 17 VDD P l=0.18u w=0.6u 
MM25 4 8 VDD VDD P l=0.18u w=0.76u 
MM24 8 CP VDD VDD P l=0.18u w=0.97u 
MM23 VDD SD 9 VDD P l=0.18u w=0.52u 
MM22 13 SC VDD VDD P l=0.18u w=0.52u 
MM21 VSS IPS QN VSS N l=0.18u w=1.03u 
MM20 17 8 IPM VSS N l=0.18u w=0.44u 
MM19 21 8 IPS VSS N l=0.18u w=0.6u 
MM17 21 3 VSS VSS N l=0.18u w=0.6u 
MM16 IPM 4 19 VSS N l=0.18u w=0.44u 
MM15 2 4 IPS VSS N l=0.18u w=0.6u 
MM14 2 IPM VSS VSS N l=0.18u w=0.75u 
MM12 24 CDN 19 VSS N l=0.18u w=0.75u 
MM18 VSS 2 24 VSS N l=0.18u w=0.75u 
MM11 3 CDN 25 VSS N l=0.18u w=1.21u 
MM13 VSS IPS 25 VSS N l=0.18u w=1.21u 
MM10 10 9 VSS VSS N l=0.18u w=0.48u 
MM9 22 10 VSS VSS N l=0.18u w=0.48u 
MM8 22 11 17 VSS N l=0.18u w=0.48u 
MM6 VSS 13 11 VSS N l=0.18u w=0.43u 
MM5 17 13 23 VSS N l=0.18u w=0.48u 
MM7 VSS D 23 VSS N l=0.18u w=0.48u 
MM2 VSS SD 9 VSS N l=0.18u w=0.43u 
MM4 4 8 VSS VSS N l=0.18u w=0.52u 
MM3 VSS CP 8 VSS N l=0.18u w=0.52u 
MM1 13 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdcrn1

.SUBCKT sdcrn2 QN  CDN CP D SC SD VDD VSS
MM43 IPM 2 19 VDD P l=0.18u w=0.6u 
MM42 IPM 3 17 VDD P l=0.18u w=0.6u 
MM41 VDD 4 19 VDD P l=0.18u w=0.55u 
MM34 19 CDN VDD VDD P l=0.18u w=0.52u 
MM40 VDD 5 21 VDD P l=0.18u w=0.76u 
MM39 IPS 3 21 VDD P l=0.18u w=0.88u 
MM37 QN IPS VDD VDD P l=0.185235u w=1.49u 
MM36 VDD IPS QN VDD P l=0.184615u w=1.482u 
MM35 VDD IPS 5 VDD P l=0.186387u w=1.146u 
MM33 VDD CDN 5 VDD P l=0.18u w=1.08u 
MM32 4 2 IPS VDD P l=0.18u w=0.88u 
MM38 4 IPM VDD VDD P l=0.18u w=0.88u 
MM31 VDD 9 10 VDD P l=0.18u w=0.52u 
MM30 22 10 VDD VDD P l=0.18u w=0.52u 
MM27 22 13 17 VDD P l=0.18u w=0.52u 
MM29 23 11 17 VDD P l=0.18u w=0.52u 
MM28 VDD D 23 VDD P l=0.18u w=0.52u 
MM26 VDD 13 11 VDD P l=0.18u w=0.5u 
MM25 3 2 VDD VDD P l=0.18u w=0.76u 
MM24 2 CP VDD VDD P l=0.18u w=0.97u 
MM23 VDD SD 9 VDD P l=0.18u w=0.52u 
MM22 13 SC VDD VDD P l=0.18u w=0.52u 
MM21 17 2 IPM VSS N l=0.18u w=0.44u 
MM20 21 2 IPS VSS N l=0.18u w=0.6u 
MM18 21 5 VSS VSS N l=0.18u w=0.6u 
MM17 IPM 3 19 VSS N l=0.18u w=0.44u 
MM16 4 3 IPS VSS N l=0.18u w=0.6u 
MM15 4 IPM VSS VSS N l=0.18u w=0.75u 
MM13 24 CDN 19 VSS N l=0.18u w=0.75u 
MM19 VSS 4 24 VSS N l=0.18u w=0.75u 
MM12 5 CDN 25 VSS N l=0.18u w=1.21u 
MM14 VSS IPS 25 VSS N l=0.18u w=1.21u 
MM11 VSS IPS QN VSS N l=0.195964u w=1.883u 
MM10 10 9 VSS VSS N l=0.18u w=0.48u 
MM9 22 10 VSS VSS N l=0.18u w=0.48u 
MM8 22 11 17 VSS N l=0.18u w=0.48u 
MM6 VSS 13 11 VSS N l=0.18u w=0.43u 
MM5 17 13 23 VSS N l=0.18u w=0.48u 
MM7 VSS D 23 VSS N l=0.18u w=0.48u 
MM2 VSS SD 9 VSS N l=0.18u w=0.43u 
MM4 3 2 VSS VSS N l=0.18u w=0.52u 
MM3 VSS CP 2 VSS N l=0.18u w=0.52u 
MM1 13 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdcrn2

.SUBCKT sdcrq1 Q  CDN CP D SC SD VDD VSS
MM42 VDD 2 19 VDD P l=0.18u w=0.55u 
MM36 19 CDN VDD VDD P l=0.18u w=0.52u 
MM41 VDD 3 20 VDD P l=0.18u w=0.76u 
MM40 IPS 4 20 VDD P l=0.18u w=0.88u 
MM37 VDD 3 Q VDD P l=0.184379u w=1.562u 
MM38 VDD IPS 3 VDD P l=0.186387u w=1.146u 
MM35 VDD CDN 3 VDD P l=0.18u w=1.08u 
MM34 2 8 IPS VDD P l=0.18u w=0.88u 
MM39 2 IPM VDD VDD P l=0.18u w=0.88u 
MM33 VDD 9 10 VDD P l=0.18u w=0.52u 
MM32 22 10 VDD VDD P l=0.18u w=0.52u 
MM29 22 13 17 VDD P l=0.18u w=0.52u 
MM31 23 11 17 VDD P l=0.18u w=0.52u 
MM30 VDD D 23 VDD P l=0.18u w=0.52u 
MM28 VDD 13 11 VDD P l=0.18u w=0.5u 
MM27 IPM 8 19 VDD P l=0.18u w=0.6u 
MM26 IPM 4 17 VDD P l=0.18u w=0.6u 
MM25 4 8 VDD VDD P l=0.18u w=0.76u 
MM24 8 CP VDD VDD P l=0.18u w=0.97u 
MM23 VDD SD 9 VDD P l=0.18u w=0.52u 
MM22 13 SC VDD VDD P l=0.18u w=0.52u 
MM21 VSS 3 Q VSS N l=0.18u w=0.98u 
MM20 17 8 IPM VSS N l=0.18u w=0.44u 
MM19 20 8 IPS VSS N l=0.18u w=0.6u 
MM17 20 3 VSS VSS N l=0.18u w=0.6u 
MM16 IPM 4 19 VSS N l=0.18u w=0.44u 
MM15 2 4 IPS VSS N l=0.18u w=0.6u 
MM14 2 IPM VSS VSS N l=0.18u w=0.75u 
MM12 24 CDN 19 VSS N l=0.18u w=0.75u 
MM18 VSS 2 24 VSS N l=0.18u w=0.75u 
MM11 3 CDN 25 VSS N l=0.18u w=1.21u 
MM13 VSS IPS 25 VSS N l=0.18u w=1.21u 
MM10 10 9 VSS VSS N l=0.18u w=0.48u 
MM9 22 10 VSS VSS N l=0.18u w=0.48u 
MM8 22 11 17 VSS N l=0.18u w=0.48u 
MM6 VSS 13 11 VSS N l=0.18u w=0.43u 
MM5 17 13 23 VSS N l=0.18u w=0.48u 
MM7 VSS D 23 VSS N l=0.18u w=0.48u 
MM2 VSS SD 9 VSS N l=0.18u w=0.43u 
MM4 4 8 VSS VSS N l=0.18u w=0.52u 
MM3 VSS CP 8 VSS N l=0.18u w=0.52u 
MM1 13 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdcrq1

.SUBCKT sdcrq2 Q  CDN CP D SC SD VDD VSS
MM43 IPM 2 19 VDD P l=0.18u w=0.6u 
MM42 IPM 3 17 VDD P l=0.18u w=0.6u 
MM41 VDD 4 19 VDD P l=0.18u w=0.55u 
MM34 19 CDN VDD VDD P l=0.18u w=0.52u 
MM40 VDD 5 21 VDD P l=0.18u w=0.76u 
MM39 IPS 3 21 VDD P l=0.18u w=0.88u 
MM36 Q 5 VDD VDD P l=0.185235u w=1.49u 
MM35 VDD 5 Q VDD P l=0.184615u w=1.482u 
MM37 VDD IPS 5 VDD P l=0.186387u w=1.146u 
MM33 VDD CDN 5 VDD P l=0.18u w=1.08u 
MM32 4 2 IPS VDD P l=0.18u w=0.88u 
MM38 4 IPM VDD VDD P l=0.18u w=0.88u 
MM31 VDD 9 10 VDD P l=0.18u w=0.52u 
MM30 22 10 VDD VDD P l=0.18u w=0.52u 
MM27 22 13 17 VDD P l=0.18u w=0.52u 
MM29 23 11 17 VDD P l=0.18u w=0.52u 
MM28 VDD D 23 VDD P l=0.18u w=0.52u 
MM26 VDD 13 11 VDD P l=0.18u w=0.5u 
MM25 3 2 VDD VDD P l=0.18u w=0.76u 
MM24 2 CP VDD VDD P l=0.18u w=0.97u 
MM23 VDD SD 9 VDD P l=0.18u w=0.52u 
MM22 13 SC VDD VDD P l=0.18u w=0.65u 
MM21 17 2 IPM VSS N l=0.18u w=0.44u 
MM20 21 2 IPS VSS N l=0.18u w=0.6u 
MM18 21 5 VSS VSS N l=0.18u w=0.6u 
MM17 IPM 3 19 VSS N l=0.18u w=0.44u 
MM16 4 3 IPS VSS N l=0.18u w=0.6u 
MM15 4 IPM VSS VSS N l=0.18u w=0.75u 
MM13 24 CDN 19 VSS N l=0.18u w=0.75u 
MM19 VSS 4 24 VSS N l=0.18u w=0.75u 
MM12 5 CDN 25 VSS N l=0.18u w=1.21u 
MM14 VSS IPS 25 VSS N l=0.18u w=1.21u 
MM11 VSS 5 Q VSS N l=0.195964u w=1.883u 
MM10 10 9 VSS VSS N l=0.18u w=0.48u 
MM9 22 10 VSS VSS N l=0.18u w=0.48u 
MM8 22 11 17 VSS N l=0.18u w=0.48u 
MM6 VSS 13 11 VSS N l=0.18u w=0.43u 
MM5 17 13 23 VSS N l=0.18u w=0.48u 
MM7 VSS D 23 VSS N l=0.18u w=0.48u 
MM2 VSS SD 9 VSS N l=0.18u w=0.43u 
MM4 3 2 VSS VSS N l=0.18u w=0.52u 
MM3 VSS CP 2 VSS N l=0.18u w=0.52u 
MM1 13 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdcrq2

.SUBCKT sdnrb1 Q QN  CP D SC SD VDD VSS
MM40 IPM 2 20 VDD P l=0.18u w=0.6u 
MM39 VDD 3 20 VDD P l=0.18u w=0.6u 
MM37 IPM 5 16 VDD P l=0.18u w=0.6u 
MM38 VDD 4 21 VDD P l=0.18u w=0.75u 
MM36 IPS 5 21 VDD P l=0.18u w=0.75u 
MM35 VDD IPM 3 VDD P l=0.18u w=0.96u 
MM33 IPS 2 3 VDD P l=0.18u w=0.84u 
MM34 4 IPS VDD VDD P l=0.186278u w=1.166u 
MM32 VDD 8 9 VDD P l=0.18u w=0.52u 
MM31 22 9 VDD VDD P l=0.18u w=0.52u 
MM28 22 12 16 VDD P l=0.18u w=0.52u 
MM30 23 10 16 VDD P l=0.18u w=0.52u 
MM29 VDD D 23 VDD P l=0.18u w=0.52u 
MM27 VDD 12 10 VDD P l=0.18u w=0.5u 
MM26 VDD 4 Q VDD P l=0.183972u w=1.722u 
MM25 VDD IPS QN VDD P l=0.183972u w=1.722u 
MM24 5 2 VDD VDD P l=0.18u w=0.76u 
MM23 2 CP VDD VDD P l=0.18u w=0.97u 
MM22 VDD SD 8 VDD P l=0.18u w=0.52u 
MM21 12 SC VDD VDD P l=0.18u w=0.7u 
MM20 16 2 IPM VSS N l=0.18u w=0.44u 
MM19 IPS 2 21 VSS N l=0.18u w=0.6u 
MM17 21 4 VSS VSS N l=0.18u w=0.6u 
MM18 VSS 3 20 VSS N l=0.18u w=0.44u 
MM16 IPM 5 20 VSS N l=0.18u w=0.44u 
MM15 3 5 IPS VSS N l=0.18u w=0.6u 
MM14 3 IPM VSS VSS N l=0.18u w=0.75u 
MM13 4 IPS VSS VSS N l=0.18u w=0.91u 
MM12 9 8 VSS VSS N l=0.18u w=0.48u 
MM11 22 9 VSS VSS N l=0.18u w=0.48u 
MM10 22 10 16 VSS N l=0.18u w=0.48u 
MM8 VSS 12 10 VSS N l=0.18u w=0.43u 
MM7 16 12 23 VSS N l=0.18u w=0.48u 
MM9 VSS D 23 VSS N l=0.18u w=0.48u 
MM4 VSS SD 8 VSS N l=0.18u w=0.43u 
MM6 5 2 VSS VSS N l=0.18u w=0.52u 
MM5 VSS CP 2 VSS N l=0.18u w=0.52u 
MM3 VSS 4 Q VSS N l=0.184743u w=1.442u 
MM2 VSS IPS QN VSS N l=0.184743u w=1.442u 
MM1 12 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdnrb1

.SUBCKT sdnrb2 Q QN  CP D SC SD VDD VSS
MM44 IPM 2 22 VDD P l=0.18u w=0.6u 
MM42 IPM 3 19 VDD P l=0.18u w=0.6u 
MM41 VDD 4 19 VDD P l=0.18u w=0.55u 
MM43 IPS 2 20 VDD P l=0.18u w=0.75u 
MM40 VDD 5 20 VDD P l=0.18u w=0.75u 
MM39 VDD IPM 4 VDD P l=0.18u w=0.96u 
MM37 IPS 3 4 VDD P l=0.18u w=0.84u 
MM38 5 IPS VDD VDD P l=0.186278u w=1.166u 
MM36 QN IPS VDD VDD P l=0.183972u w=1.722u 
MM35 QN IPS VDD VDD P l=0.183972u w=1.722u 
MM34 Q 5 VDD VDD P l=0.183972u w=1.722u 
MM33 VDD 5 Q VDD P l=0.183972u w=1.722u 
MM32 VDD 8 9 VDD P l=0.18u w=0.52u 
MM31 21 9 VDD VDD P l=0.18u w=0.52u 
MM28 21 12 22 VDD P l=0.18u w=0.52u 
MM30 23 10 22 VDD P l=0.18u w=0.52u 
MM29 VDD D 23 VDD P l=0.18u w=0.52u 
MM27 VDD 12 10 VDD P l=0.18u w=0.5u 
MM26 2 3 VDD VDD P l=0.18u w=0.76u 
MM25 3 CP VDD VDD P l=0.18u w=0.97u 
MM24 VDD SD 8 VDD P l=0.18u w=0.52u 
MM23 12 SC VDD VDD P l=0.18u w=0.52u 
MM22 IPM 2 19 VSS N l=0.18u w=0.44u 
MM20 22 3 IPM VSS N l=0.18u w=0.44u 
MM21 4 2 IPS VSS N l=0.18u w=0.6u 
MM19 IPS 3 20 VSS N l=0.18u w=0.6u 
MM18 VSS 4 19 VSS N l=0.18u w=0.44u 
MM17 20 5 VSS VSS N l=0.18u w=0.6u 
MM16 4 IPM VSS VSS N l=0.18u w=0.75u 
MM15 5 IPS VSS VSS N l=0.18u w=0.91u 
MM14 QN IPS VSS VSS N l=0.184743u w=1.442u 
MM13 QN IPS VSS VSS N l=0.184743u w=1.442u 
MM12 VSS 5 Q VSS N l=0.184743u w=1.442u 
MM11 Q 5 VSS VSS N l=0.184743u w=1.442u 
MM10 9 8 VSS VSS N l=0.18u w=0.48u 
MM9 21 9 VSS VSS N l=0.18u w=0.48u 
MM8 21 10 22 VSS N l=0.18u w=0.48u 
MM6 VSS 12 10 VSS N l=0.18u w=0.43u 
MM5 22 12 23 VSS N l=0.18u w=0.48u 
MM7 VSS D 23 VSS N l=0.18u w=0.48u 
MM2 VSS SD 8 VSS N l=0.18u w=0.43u 
MM4 2 3 VSS VSS N l=0.18u w=0.52u 
MM3 VSS CP 3 VSS N l=0.18u w=0.52u 
MM1 12 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdnrb2

.SUBCKT sdnrn1 QN  CP D SC SD VDD VSS
MM38 6 2 VDD VDD P l=0.18u w=0.76u 
MM37 2 CP VDD VDD P l=0.18u w=0.97u 
MM36 IPM 2 19 VDD P l=0.18u w=0.6u 
MM35 VDD 4 19 VDD P l=0.18u w=0.55u 
MM33 IPM 6 16 VDD P l=0.18u w=0.6u 
MM34 VDD 5 20 VDD P l=0.18u w=0.75u 
MM32 IPS 6 20 VDD P l=0.18u w=0.75u 
MM31 VDD IPM 4 VDD P l=0.18u w=0.96u 
MM29 IPS 2 4 VDD P l=0.18u w=0.84u 
MM30 VDD IPS 5 VDD P l=0.18u w=0.75u 
MM28 VDD 9 10 VDD P l=0.18u w=0.52u 
MM27 21 10 VDD VDD P l=0.18u w=0.52u 
MM24 21 13 16 VDD P l=0.18u w=0.52u 
MM26 22 11 16 VDD P l=0.18u w=0.52u 
MM25 VDD D 22 VDD P l=0.18u w=0.52u 
MM23 VDD 13 11 VDD P l=0.18u w=0.5u 
MM22 QN IPS VDD VDD P l=0.184217u w=1.622u 
MM21 VDD SD 9 VDD P l=0.18u w=0.52u 
MM20 13 SC VDD VDD P l=0.18u w=0.52u 
MM17 VSS SD 9 VSS N l=0.18u w=0.43u 
MM19 6 2 VSS VSS N l=0.18u w=0.52u 
MM18 VSS CP 2 VSS N l=0.18u w=0.52u 
MM16 16 2 IPM VSS N l=0.18u w=0.44u 
MM15 IPS 2 20 VSS N l=0.18u w=0.6u 
MM13 20 5 VSS VSS N l=0.18u w=0.6u 
MM14 VSS 4 19 VSS N l=0.18u w=0.44u 
MM12 IPM 6 19 VSS N l=0.18u w=0.44u 
MM11 4 6 IPS VSS N l=0.18u w=0.6u 
MM10 4 IPM VSS VSS N l=0.18u w=0.75u 
MM9 5 IPS VSS VSS N l=0.18u w=0.6u 
MM8 10 9 VSS VSS N l=0.18u w=0.48u 
MM7 21 10 VSS VSS N l=0.18u w=0.48u 
MM6 21 11 16 VSS N l=0.18u w=0.48u 
MM4 VSS 13 11 VSS N l=0.18u w=0.43u 
MM3 16 13 22 VSS N l=0.18u w=0.48u 
MM5 VSS D 22 VSS N l=0.18u w=0.48u 
MM2 QN IPS VSS VSS N l=0.185886u w=1.162u 
MM1 13 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdnrn1

.SUBCKT sdnrn2 QN  CP D SC SD VDD VSS
MM40 IPM 2 19 VDD P l=0.18u w=0.6u 
MM39 VDD 3 19 VDD P l=0.18u w=0.55u 
MM37 IPM 5 16 VDD P l=0.18u w=0.6u 
MM38 VDD 4 20 VDD P l=0.18u w=0.75u 
MM36 IPS 5 20 VDD P l=0.18u w=0.75u 
MM35 VDD IPM 3 VDD P l=0.18u w=0.96u 
MM33 IPS 2 3 VDD P l=0.18u w=0.84u 
MM34 4 IPS VDD VDD P l=0.186278u w=1.166u 
MM32 VDD 8 9 VDD P l=0.18u w=0.52u 
MM31 21 9 VDD VDD P l=0.18u w=0.52u 
MM28 21 12 16 VDD P l=0.18u w=0.52u 
MM30 22 10 16 VDD P l=0.18u w=0.52u 
MM29 VDD D 22 VDD P l=0.18u w=0.52u 
MM27 VDD 12 10 VDD P l=0.18u w=0.5u 
MM26 QN IPS VDD VDD P l=0.183972u w=1.722u 
MM25 QN IPS VDD VDD P l=0.184241u w=1.726u 
MM24 5 2 VDD VDD P l=0.18u w=0.76u 
MM23 2 CP VDD VDD P l=0.18u w=0.97u 
MM22 VDD SD 8 VDD P l=0.18u w=0.52u 
MM21 12 SC VDD VDD P l=0.18u w=0.52u 
MM20 QN IPS VSS VSS N l=0.184743u w=1.442u 
MM19 QN IPS VSS VSS N l=0.184743u w=1.442u 
MM18 16 2 IPM VSS N l=0.18u w=0.44u 
MM17 IPS 2 20 VSS N l=0.18u w=0.6u 
MM15 20 4 VSS VSS N l=0.18u w=0.6u 
MM16 VSS 3 19 VSS N l=0.18u w=0.44u 
MM14 IPM 5 19 VSS N l=0.18u w=0.44u 
MM13 3 5 IPS VSS N l=0.18u w=0.6u 
MM12 3 IPM VSS VSS N l=0.18u w=0.75u 
MM11 4 IPS VSS VSS N l=0.18u w=0.91u 
MM10 9 8 VSS VSS N l=0.18u w=0.48u 
MM9 21 9 VSS VSS N l=0.18u w=0.48u 
MM8 21 10 16 VSS N l=0.18u w=0.48u 
MM6 VSS 12 10 VSS N l=0.18u w=0.43u 
MM5 16 12 22 VSS N l=0.18u w=0.48u 
MM7 VSS D 22 VSS N l=0.18u w=0.48u 
MM2 VSS SD 8 VSS N l=0.18u w=0.43u 
MM4 5 2 VSS VSS N l=0.18u w=0.52u 
MM3 VSS CP 2 VSS N l=0.18u w=0.52u 
MM1 12 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdnrn2

.SUBCKT sdnrq1 Q  CP D SC SD VDD VSS
MM38 VDD 2 7 VDD P l=0.18u w=0.81u 
MM37 VDD CP 2 VDD P l=0.186618u w=1.106u 
MM36 4 2 15 VDD P l=0.18u w=0.78u 
MM30 15 7 20 VDD P l=0.18u w=0.57u 
MM35 IPM 2 19 VDD P l=0.18u w=0.42u 
MM34 VDD 4 19 VDD P l=0.18u w=0.42u 
MM32 4 IPM VDD VDD P l=0.18u w=0.78u 
MM31 16 7 IPM VDD P l=0.18u w=0.51u 
MM33 VDD IPS 20 VDD P l=0.18u w=0.5u 
MM29 13 SC VDD VDD P l=0.18u w=0.5u 
MM28 10 9 VDD VDD P l=0.18u w=0.51u 
MM27 21 10 VDD VDD P l=0.18u w=0.51u 
MM24 21 13 16 VDD P l=0.18u w=0.59u 
MM26 VDD D 22 VDD P l=0.18u w=0.59u 
MM25 16 12 22 VDD P l=0.18u w=0.59u 
MM23 VDD 13 12 VDD P l=0.18u w=0.5u 
MM22 9 SD VDD VDD P l=0.18u w=0.5u 
MM21 VDD 15 IPS VDD P l=0.18u w=1.05u 
MM20 Q IPS VDD VDD P l=0.184586u w=1.596u 
MM19 7 2 VSS VSS N l=0.18u w=0.5u 
MM18 VSS CP 2 VSS N l=0.18u w=0.5u 
MM17 16 2 IPM VSS N l=0.18u w=0.84u 
MM16 15 2 20 VSS N l=0.18u w=0.77u 
MM14 VSS IPS 20 VSS N l=0.18u w=0.77u 
MM15 VSS 4 19 VSS N l=0.18u w=0.84u 
MM12 19 7 IPM VSS N l=0.18u w=0.84u 
MM11 VSS 15 IPS VSS N l=0.18u w=0.77u 
MM10 4 7 15 VSS N l=0.18u w=0.77u 
MM13 4 IPM VSS VSS N l=0.18u w=0.77u 
MM9 VSS SD 9 VSS N l=0.18u w=0.42u 
MM8 10 9 VSS VSS N l=0.18u w=0.48u 
MM7 21 10 VSS VSS N l=0.18u w=0.84u 
MM5 21 12 16 VSS N l=0.18u w=0.84u 
MM4 12 13 VSS VSS N l=0.18u w=0.48u 
MM3 22 13 16 VSS N l=0.18u w=0.84u 
MM6 22 D VSS VSS N l=0.18u w=0.84u 
MM2 Q IPS VSS VSS N l=0.18u w=1.2u 
MM1 13 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdnrq1

.SUBCKT sdnrq2 Q  CP D SC SD VDD VSS
MM40 VDD 2 7 VDD P l=0.18u w=0.81u 
MM39 VDD CP 2 VDD P l=0.186618u w=1.106u 
MM38 4 2 15 VDD P l=0.18u w=0.78u 
MM32 15 7 20 VDD P l=0.18u w=0.57u 
MM37 IPM 2 19 VDD P l=0.18u w=0.42u 
MM36 VDD 4 19 VDD P l=0.18u w=0.42u 
MM34 4 IPM VDD VDD P l=0.18u w=0.78u 
MM33 16 7 IPM VDD P l=0.18u w=0.51u 
MM35 VDD IPS 20 VDD P l=0.18u w=0.5u 
MM31 13 SC VDD VDD P l=0.18u w=0.5u 
MM30 10 9 VDD VDD P l=0.18u w=0.51u 
MM29 21 10 VDD VDD P l=0.18u w=0.51u 
MM26 21 13 16 VDD P l=0.18u w=0.59u 
MM28 VDD D 22 VDD P l=0.18u w=0.59u 
MM27 16 12 22 VDD P l=0.18u w=0.59u 
MM25 VDD 13 12 VDD P l=0.18u w=0.5u 
MM24 9 SD VDD VDD P l=0.18u w=0.5u 
MM23 VDD 15 IPS VDD P l=0.186964u w=1.12u 
MM22 Q IPS VDD VDD P l=0.185162u w=1.604u 
MM21 Q IPS VDD VDD P l=0.18u w=1.53u 
MM20 7 2 VSS VSS N l=0.18u w=0.5u 
MM19 VSS CP 2 VSS N l=0.18u w=0.5u 
MM18 16 2 IPM VSS N l=0.18u w=0.84u 
MM17 15 2 20 VSS N l=0.18u w=0.77u 
MM15 VSS IPS 20 VSS N l=0.18u w=0.77u 
MM16 VSS 4 19 VSS N l=0.18u w=0.84u 
MM13 19 7 IPM VSS N l=0.18u w=0.84u 
MM12 VSS 15 IPS VSS N l=0.18u w=0.77u 
MM11 4 7 15 VSS N l=0.18u w=0.77u 
MM14 4 IPM VSS VSS N l=0.18u w=0.77u 
MM10 VSS SD 9 VSS N l=0.18u w=0.42u 
MM9 10 9 VSS VSS N l=0.18u w=0.48u 
MM8 21 10 VSS VSS N l=0.18u w=0.84u 
MM6 21 12 16 VSS N l=0.18u w=0.84u 
MM5 12 13 VSS VSS N l=0.18u w=0.48u 
MM4 22 13 16 VSS N l=0.18u w=0.84u 
MM7 22 D VSS VSS N l=0.18u w=0.84u 
MM3 Q IPS VSS VSS N l=0.186499u w=1.274u 
MM2 Q IPS VSS VSS N l=0.18u w=1.2u 
MM1 13 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdnrq2

.SUBCKT sdprb1 Q QN  CP D SC SD SDN VDD VSS
MM44 23 2 IPM VDD P l=0.18u w=0.51u 
MM43 IPM 3 18 VDD P l=0.18u w=0.51u 
MM42 VDD 4 18 VDD P l=0.18u w=0.51u 
MM41 VDD 3 2 VDD P l=0.18u w=0.81u 
MM40 VDD CP 3 VDD P l=0.186618u w=1.106u 
MM39 11 SC VDD VDD P l=0.18u w=0.5u 
MM38 8 7 VDD VDD P l=0.18u w=0.51u 
MM37 22 8 VDD VDD P l=0.18u w=0.51u 
MM34 22 11 23 VDD P l=0.18u w=0.59u 
MM36 VDD D 24 VDD P l=0.18u w=0.59u 
MM35 23 10 24 VDD P l=0.18u w=0.59u 
MM33 VDD 11 10 VDD P l=0.18u w=0.5u 
MM32 7 SD VDD VDD P l=0.18u w=0.5u 
MM31 VDD 13 Q VDD P l=0.18u w=1.5u 
MM30 13 IPS VDD VDD P l=0.185971u w=1.226u 
MM29 QN IPS VDD VDD P l=0.18u w=1.5u 
MM28 21 2 IPS VDD P l=0.18u w=0.78u 
MM25 21 SDN VDD VDD P l=0.186042u w=1.132u 
MM27 4 IPM VDD VDD P l=0.186502u w=1.052u 
MM26 21 13 VDD VDD P l=0.186042u w=1.132u 
MM24 4 SDN VDD VDD P l=0.186502u w=1.052u 
MM23 4 3 IPS VDD P l=0.18u w=0.78u 
MM20 23 3 IPM VSS N l=0.18u w=0.76u 
MM22 18 2 IPM VSS N l=0.18u w=0.76u 
MM21 4 2 IPS VSS N l=0.18u w=0.76u 
MM19 21 3 IPS VSS N l=0.18u w=0.76u 
MM18 VSS 4 18 VSS N l=0.18u w=0.76u 
MM15 21 SDN 25 VSS N l=0.18u w=0.95u 
MM16 VSS 13 25 VSS N l=0.18u w=0.95u 
MM14 26 SDN 4 VSS N l=0.18u w=0.95u 
MM17 26 IPM VSS VSS N l=0.18u w=0.95u 
MM13 VSS IPS 13 VSS N l=0.18u w=0.95u 
MM12 VSS 13 Q VSS N l=0.18u w=1.08u 
MM11 VSS IPS QN VSS N l=0.18u w=1.08u 
MM10 VSS SD 7 VSS N l=0.18u w=0.42u 
MM9 8 7 VSS VSS N l=0.18u w=0.48u 
MM8 22 8 VSS VSS N l=0.18u w=0.84u 
MM6 22 10 23 VSS N l=0.18u w=0.84u 
MM5 10 11 VSS VSS N l=0.18u w=0.48u 
MM4 24 11 23 VSS N l=0.18u w=0.84u 
MM7 24 D VSS VSS N l=0.18u w=0.84u 
MM3 2 3 VSS VSS N l=0.18u w=0.5u 
MM2 VSS CP 3 VSS N l=0.18u w=0.5u 
MM1 11 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdprb1

.SUBCKT sdprb2 Q QN  CP D SC SD SDN VDD VSS
MM48 23 2 IPM VDD P l=0.18u w=0.51u 
MM47 IPM 3 17 VDD P l=0.18u w=0.51u 
MM46 VDD 4 17 VDD P l=0.18u w=0.51u 
MM45 VDD 5 Q VDD P l=0.18u w=1.5u 
MM44 Q 5 VDD VDD P l=0.18u w=1.5u 
MM43 5 IPS VDD VDD P l=0.185971u w=1.226u 
MM42 VDD IPS QN VDD P l=0.18u w=1.5u 
MM41 QN IPS VDD VDD P l=0.18u w=1.5u 
MM40 VDD 3 2 VDD P l=0.18u w=0.81u 
MM39 VDD CP 3 VDD P l=0.186618u w=1.106u 
MM38 13 SC VDD VDD P l=0.18u w=0.5u 
MM37 10 9 VDD VDD P l=0.18u w=0.51u 
MM36 22 10 VDD VDD P l=0.18u w=0.51u 
MM33 22 13 23 VDD P l=0.18u w=0.59u 
MM35 VDD D 24 VDD P l=0.18u w=0.59u 
MM34 23 12 24 VDD P l=0.18u w=0.59u 
MM32 VDD 13 12 VDD P l=0.18u w=0.5u 
MM31 9 SD VDD VDD P l=0.18u w=0.5u 
MM30 21 2 IPS VDD P l=0.18u w=0.78u 
MM27 21 SDN VDD VDD P l=0.186042u w=1.132u 
MM29 4 IPM VDD VDD P l=0.186502u w=1.052u 
MM28 21 5 VDD VDD P l=0.186042u w=1.132u 
MM26 4 SDN VDD VDD P l=0.186502u w=1.052u 
MM25 4 3 IPS VDD P l=0.18u w=0.78u 
MM22 23 3 IPM VSS N l=0.18u w=0.76u 
MM24 17 2 IPM VSS N l=0.18u w=0.76u 
MM23 4 2 IPS VSS N l=0.18u w=0.76u 
MM21 21 3 IPS VSS N l=0.18u w=0.76u 
MM20 VSS 4 17 VSS N l=0.18u w=0.76u 
MM17 21 SDN 25 VSS N l=0.18u w=0.95u 
MM18 VSS 5 25 VSS N l=0.18u w=0.95u 
MM16 26 SDN 4 VSS N l=0.18u w=0.95u 
MM19 26 IPM VSS VSS N l=0.18u w=0.95u 
MM15 VSS IPS 5 VSS N l=0.18u w=0.95u 
MM14 VSS 5 Q VSS N l=0.18u w=1.08u 
MM13 VSS 5 Q VSS N l=0.18u w=1.08u 
MM12 QN IPS VSS VSS N l=0.18u w=1.08u 
MM11 QN IPS VSS VSS N l=0.18u w=1.08u 
MM10 VSS SD 9 VSS N l=0.18u w=0.42u 
MM9 10 9 VSS VSS N l=0.18u w=0.48u 
MM8 22 10 VSS VSS N l=0.18u w=0.84u 
MM6 22 12 23 VSS N l=0.18u w=0.84u 
MM5 12 13 VSS VSS N l=0.18u w=0.48u 
MM4 24 13 23 VSS N l=0.18u w=0.84u 
MM7 24 D VSS VSS N l=0.18u w=0.84u 
MM3 2 3 VSS VSS N l=0.18u w=0.5u 
MM2 VSS CP 3 VSS N l=0.18u w=0.5u 
MM1 13 SC VSS VSS N l=0.18u w=0.48u 
.ENDS sdprb2

.SUBCKT secrq1 Q  CDN CP D ENN SC SD VDD VSS
MM59 VDD D 29 VDD P l=0.18u w=0.64u 
MM58 24 4 29 VDD P l=0.18u w=0.58u 
MM49 VDD IPS 6 VDD P l=0.18u w=1.23u 
MM48 6 CDN VDD VDD P l=0.18635u w=1.304u 
MM41 14 15 VDD VDD P l=0.18u w=0.98u 
MM33 VDD SC 16 VDD P l=0.18u w=0.6u 
MM32 VDD SD 15 VDD P l=0.18u w=0.86u 
MM31 VDD 16 22 VDD P l=0.18u w=0.64u 
MM40 24 16 30 VDD P l=0.18u w=0.52u 
MM42 VDD 14 30 VDD P l=0.18u w=0.52u 
MM39 VDD ENN 18 VDD P l=0.18u w=0.52u 
MM37 2 ENN VDD VDD P l=0.186783u w=1.15u 
MM35 VDD 16 2 VDD P l=0.186387u w=1.146u 
MM57 24 2 25 VDD P l=0.18u w=0.58u 
MM36 VDD 4 23 VDD P l=0.18u w=0.52u 
MM38 VDD 18 4 VDD P l=0.18u w=0.52u 
MM34 VDD 16 4 VDD P l=0.18u w=0.52u 
MM60 VDD 2 21 VDD P l=0.18u w=0.52u 
MM45 VDD CP 9 VDD P l=0.187156u w=1.09u 
MM43 25 13 VDD VDD P l=0.18u w=0.57u 
MM56 28 5 VDD VDD P l=0.187631u w=1.148u 
MM53 24 8 IPM VDD P l=0.18u w=0.54u 
MM51 28 9 IPM VDD P l=0.18u w=0.54u 
MM47 28 CDN VDD VDD P l=0.18u w=0.98u 
MM44 VDD 9 8 VDD P l=0.18u w=1.02u 
MM55 VDD 6 13 VDD P l=0.18u w=0.67u 
MM52 IPS 8 13 VDD P l=0.18u w=0.67u 
MM46 IPS 9 5 VDD P l=0.18u w=0.67u 
MM54 5 IPM VDD VDD P l=0.18u w=0.67u 
MM50 VDD 6 Q VDD P l=0.18u w=1.5u 
MM21 5 8 IPS VSS N l=0.18u w=0.49u 
MM19 13 9 IPS VSS N l=0.18u w=0.49u 
MM12 VSS ENN 18 VSS N l=0.18u w=0.44u 
MM9 2 ENN 32 VSS N l=0.18u w=0.49u 
MM6 24 22 30 VSS N l=0.18u w=0.44u 
MM5 VSS 14 30 VSS N l=0.18u w=0.44u 
MM4 VSS 15 14 VSS N l=0.18u w=0.96u 
MM3 VSS 16 22 VSS N l=0.18u w=0.44u 
MM2 16 SC VSS VSS N l=0.18u w=0.65u 
MM1 15 SD VSS VSS N l=0.18u w=0.64u 
MM30 25 21 24 VSS N l=0.18u w=0.44u 
MM29 21 2 VSS VSS N l=0.18u w=0.44u 
MM28 24 23 29 VSS N l=0.18u w=0.44u 
MM27 29 D VSS VSS N l=0.18u w=0.44u 
MM11 23 4 VSS VSS N l=0.18u w=0.44u 
MM10 4 18 31 VSS N l=0.18u w=0.44u 
MM8 VSS 16 31 VSS N l=0.18u w=0.44u 
MM7 VSS 16 32 VSS N l=0.18u w=0.49u 
MM26 25 13 VSS VSS N l=0.18u w=0.44u 
MM20 IPM 9 24 VSS N l=0.18u w=0.45u 
MM23 VSS IPM 5 VSS N l=0.18u w=0.57u 
MM22 28 8 IPM VSS N l=0.18u w=0.6u 
MM16 33 CDN 28 VSS N l=0.18u w=0.49u 
MM25 VSS 5 33 VSS N l=0.18u w=0.49u 
MM14 VSS CP 9 VSS N l=0.186803u w=1.076u 
MM13 VSS 9 8 VSS N l=0.18u w=0.96u 
MM24 VSS 6 13 VSS N l=0.18u w=0.57u 
MM18 VSS 6 Q VSS N l=0.18u w=1u 
MM15 34 CDN 6 VSS N l=0.18u w=0.98u 
MM17 VSS IPS 34 VSS N l=0.18u w=0.98u 
.ENDS secrq1

.SUBCKT secrq2 Q  CDN CP D ENN SC SD VDD VSS
MM61 VDD D 29 VDD P l=0.18u w=0.64u 
MM60 24 4 29 VDD P l=0.18u w=0.58u 
MM45 VDD 9 8 VDD P l=0.18u w=1.02u 
MM42 14 15 VDD VDD P l=0.18u w=0.98u 
MM34 VDD SC 16 VDD P l=0.18u w=0.6u 
MM33 VDD SD 15 VDD P l=0.18u w=0.86u 
MM32 VDD 16 22 VDD P l=0.18u w=0.64u 
MM41 24 16 30 VDD P l=0.18u w=0.52u 
MM43 VDD 14 30 VDD P l=0.18u w=0.52u 
MM40 VDD ENN 18 VDD P l=0.18u w=0.52u 
MM38 2 ENN VDD VDD P l=0.186783u w=1.15u 
MM36 VDD 16 2 VDD P l=0.186387u w=1.146u 
MM59 24 2 25 VDD P l=0.18u w=0.58u 
MM37 VDD 4 23 VDD P l=0.18u w=0.52u 
MM39 VDD 18 4 VDD P l=0.18u w=0.52u 
MM35 VDD 16 4 VDD P l=0.18u w=0.52u 
MM62 VDD 2 21 VDD P l=0.18u w=0.52u 
MM46 VDD CP 9 VDD P l=0.187156u w=1.09u 
MM44 25 13 VDD VDD P l=0.18u w=0.57u 
MM58 28 5 VDD VDD P l=0.187631u w=1.148u 
MM55 24 8 IPM VDD P l=0.18u w=0.54u 
MM53 28 9 IPM VDD P l=0.18u w=0.54u 
MM48 28 CDN VDD VDD P l=0.18u w=0.98u 
MM57 VDD 6 13 VDD P l=0.18u w=0.67u 
MM54 IPS 8 13 VDD P l=0.18u w=0.67u 
MM50 VDD IPS 6 VDD P l=0.18u w=1.23u 
MM49 6 CDN VDD VDD P l=0.18635u w=1.304u 
MM47 IPS 9 5 VDD P l=0.18u w=0.67u 
MM56 5 IPM VDD VDD P l=0.18u w=0.67u 
MM52 VDD 6 Q VDD P l=0.18526u w=1.574u 
MM51 VDD 6 Q VDD P l=0.18u w=1.5u 
MM22 5 8 IPS VSS N l=0.18u w=0.49u 
MM20 13 9 IPS VSS N l=0.18u w=0.49u 
MM12 VSS ENN 18 VSS N l=0.18u w=0.44u 
MM9 2 ENN 32 VSS N l=0.18u w=0.49u 
MM6 24 22 30 VSS N l=0.18u w=0.44u 
MM5 VSS 14 30 VSS N l=0.18u w=0.44u 
MM4 VSS 15 14 VSS N l=0.18u w=0.96u 
MM3 VSS 16 22 VSS N l=0.18u w=0.44u 
MM2 16 SC VSS VSS N l=0.18u w=0.65u 
MM1 15 SD VSS VSS N l=0.18u w=0.64u 
MM31 21 2 VSS VSS N l=0.18u w=0.44u 
MM30 25 21 24 VSS N l=0.18u w=0.44u 
MM29 24 23 29 VSS N l=0.18u w=0.44u 
MM28 29 D VSS VSS N l=0.18u w=0.44u 
MM11 23 4 VSS VSS N l=0.18u w=0.44u 
MM10 4 18 31 VSS N l=0.18u w=0.44u 
MM8 VSS 16 31 VSS N l=0.18u w=0.44u 
MM7 VSS 16 32 VSS N l=0.18u w=0.49u 
MM27 25 13 VSS VSS N l=0.18u w=0.44u 
MM21 IPM 9 24 VSS N l=0.18u w=0.45u 
MM24 VSS IPM 5 VSS N l=0.18u w=0.57u 
MM23 28 8 IPM VSS N l=0.18u w=0.6u 
MM16 33 CDN 28 VSS N l=0.18u w=0.49u 
MM26 VSS 5 33 VSS N l=0.18u w=0.49u 
MM14 VSS CP 9 VSS N l=0.186803u w=1.076u 
MM13 VSS 9 8 VSS N l=0.18u w=0.96u 
MM25 VSS 6 13 VSS N l=0.18u w=0.57u 
MM19 Q 6 VSS VSS N l=0.187113u w=1.164u 
MM18 VSS 6 Q VSS N l=0.18u w=1.09u 
MM15 34 CDN 6 VSS N l=0.18u w=0.98u 
MM17 VSS IPS 34 VSS N l=0.18u w=0.98u 
.ENDS secrq2

.SUBCKT senrq1 Q  CP D ENN SC SD VDD VSS
MM52 VDD CP 6 VDD P l=0.188434u w=1.245u 
MM38 VDD IPS 8 VDD P l=0.184171u w=1.87u 
MM41 12 13 VDD VDD P l=0.18u w=0.98u 
MM40 24 14 29 VDD P l=0.18u w=0.52u 
MM42 VDD 12 29 VDD P l=0.18u w=0.52u 
MM37 VDD ENN 17 VDD P l=0.18u w=0.52u 
MM35 3 ENN VDD VDD P l=0.186783u w=1.15u 
MM33 VDD 14 3 VDD P l=0.186387u w=1.146u 
MM31 VDD SC 14 VDD P l=0.18u w=0.6u 
MM30 VDD SD 13 VDD P l=0.18u w=0.86u 
MM29 VDD 14 21 VDD P l=0.18u w=0.64u 
MM56 VDD D 23 VDD P l=0.18u w=0.64u 
MM54 24 4 23 VDD P l=0.18u w=0.58u 
MM55 VDD 3 20 VDD P l=0.18u w=0.52u 
MM53 24 3 25 VDD P l=0.18u w=0.58u 
MM43 25 11 VDD VDD P l=0.18u w=0.57u 
MM34 VDD 4 22 VDD P l=0.18u w=0.52u 
MM36 VDD 17 4 VDD P l=0.18u w=0.52u 
MM32 VDD 14 4 VDD P l=0.18u w=0.52u 
MM51 VDD 6 10 VDD P l=0.18u w=1.26u 
MM48 7 IPM VDD VDD P l=0.18u w=0.75u 
MM45 7 6 IPS VDD P l=0.18u w=0.6u 
MM47 IPM 10 24 VDD P l=0.18u w=0.52u 
MM49 11 8 VDD VDD P l=0.18u w=0.6u 
MM46 11 10 IPS VDD P l=0.18u w=0.6u 
MM50 VDD 7 27 VDD P l=0.18u w=0.52u 
MM44 IPM 6 27 VDD P l=0.18u w=0.52u 
MM39 VDD 8 Q VDD P l=0.18u w=1.8u 
MM23 11 8 VSS VSS N l=0.18u w=0.47u 
MM18 11 6 IPS VSS N l=0.18u w=0.47u 
MM14 VSS ENN 17 VSS N l=0.18u w=0.44u 
MM11 3 ENN 31 VSS N l=0.18u w=0.49u 
MM8 24 21 29 VSS N l=0.18u w=0.44u 
MM7 VSS 12 29 VSS N l=0.18u w=0.44u 
MM6 VSS 13 12 VSS N l=0.18u w=0.96u 
MM3 VSS 14 21 VSS N l=0.18u w=0.44u 
MM2 14 SC VSS VSS N l=0.18u w=0.65u 
MM1 13 SD VSS VSS N l=0.18u w=0.64u 
MM27 25 20 24 VSS N l=0.18u w=0.44u 
MM26 20 3 VSS VSS N l=0.18u w=0.44u 
MM28 23 D VSS VSS N l=0.18u w=0.44u 
MM25 24 22 23 VSS N l=0.18u w=0.44u 
MM13 22 4 VSS VSS N l=0.18u w=0.44u 
MM12 4 17 30 VSS N l=0.18u w=0.44u 
MM10 VSS 14 30 VSS N l=0.18u w=0.44u 
MM9 VSS 14 31 VSS N l=0.18u w=0.49u 
MM19 IPM 6 24 VSS N l=0.18u w=0.52u 
MM24 27 7 VSS VSS N l=0.18u w=0.47u 
MM21 IPM 10 27 VSS N l=0.18u w=0.52u 
MM22 7 IPM VSS VSS N l=0.18u w=0.47u 
MM20 IPS 10 7 VSS N l=0.18u w=0.47u 
MM17 25 11 VSS VSS N l=0.18u w=0.44u 
MM16 VSS CP 6 VSS N l=0.187906u w=1.108u 
MM15 VSS 6 10 VSS N l=0.18u w=0.97u 
MM5 VSS 8 Q VSS N l=0.18u w=1.21u 
MM4 VSS IPS 8 VSS N l=0.186094u w=1.28u 
.ENDS senrq1

.SUBCKT senrq2 Q  CP D ENN SC SD VDD VSS
MM49 IPM 10 23 VDD P l=0.18u w=0.52u 
MM46 IPM 6 26 VDD P l=0.18u w=0.52u 
MM43 12 13 VDD VDD P l=0.18u w=0.98u 
MM42 23 14 29 VDD P l=0.18u w=0.52u 
MM44 VDD 12 29 VDD P l=0.18u w=0.52u 
MM38 VDD ENN 17 VDD P l=0.18u w=0.52u 
MM36 3 ENN VDD VDD P l=0.186783u w=1.15u 
MM34 VDD 14 3 VDD P l=0.186387u w=1.146u 
MM37 VDD 17 4 VDD P l=0.18u w=0.52u 
MM33 VDD 14 4 VDD P l=0.18u w=0.52u 
MM32 VDD SC 14 VDD P l=0.18u w=0.6u 
MM31 VDD SD 13 VDD P l=0.18u w=0.86u 
MM30 VDD 14 21 VDD P l=0.18u w=0.64u 
MM58 VDD D 28 VDD P l=0.18u w=0.64u 
MM56 23 4 28 VDD P l=0.18u w=0.58u 
MM57 VDD 3 20 VDD P l=0.18u w=0.52u 
MM55 23 3 24 VDD P l=0.18u w=0.58u 
MM54 VDD CP 6 VDD P l=0.188434u w=1.245u 
MM53 VDD 6 10 VDD P l=0.18u w=1.26u 
MM45 24 11 VDD VDD P l=0.18u w=0.57u 
MM35 VDD 4 22 VDD P l=0.18u w=0.52u 
MM50 7 IPM VDD VDD P l=0.18u w=0.75u 
MM47 7 6 IPS VDD P l=0.18u w=0.6u 
MM51 11 8 VDD VDD P l=0.18u w=0.6u 
MM48 11 10 IPS VDD P l=0.18u w=0.6u 
MM52 VDD 7 26 VDD P l=0.18u w=0.52u 
MM41 Q 8 VDD VDD P l=0.184171u w=1.87u 
MM40 VDD 8 Q VDD P l=0.18u w=1.8u 
MM39 VDD IPS 8 VDD P l=0.184171u w=1.87u 
MM24 11 8 VSS VSS N l=0.18u w=0.47u 
MM19 11 6 IPS VSS N l=0.18u w=0.47u 
MM15 VSS ENN 17 VSS N l=0.18u w=0.44u 
MM12 3 ENN 31 VSS N l=0.18u w=0.49u 
MM9 23 21 29 VSS N l=0.18u w=0.44u 
MM8 VSS 12 29 VSS N l=0.18u w=0.44u 
MM7 VSS 13 12 VSS N l=0.18u w=0.96u 
MM3 VSS 14 21 VSS N l=0.18u w=0.44u 
MM2 14 SC VSS VSS N l=0.18u w=0.65u 
MM1 13 SD VSS VSS N l=0.18u w=0.64u 
MM28 24 20 23 VSS N l=0.18u w=0.44u 
MM27 20 3 VSS VSS N l=0.18u w=0.44u 
MM29 28 D VSS VSS N l=0.18u w=0.44u 
MM26 23 22 28 VSS N l=0.18u w=0.44u 
MM14 22 4 VSS VSS N l=0.18u w=0.44u 
MM13 4 17 30 VSS N l=0.18u w=0.44u 
MM11 VSS 14 30 VSS N l=0.18u w=0.44u 
MM10 VSS 14 31 VSS N l=0.18u w=0.49u 
MM20 IPM 6 23 VSS N l=0.18u w=0.52u 
MM25 26 7 VSS VSS N l=0.18u w=0.47u 
MM22 IPM 10 26 VSS N l=0.18u w=0.52u 
MM23 7 IPM VSS VSS N l=0.18u w=0.47u 
MM21 IPS 10 7 VSS N l=0.18u w=0.47u 
MM18 24 11 VSS VSS N l=0.18u w=0.44u 
MM17 VSS CP 6 VSS N l=0.187906u w=1.108u 
MM16 VSS 6 10 VSS N l=0.18u w=0.97u 
MM6 VSS 8 Q VSS N l=0.186094u w=1.28u 
MM5 VSS 8 Q VSS N l=0.18u w=1.21u 
MM4 VSS IPS 8 VSS N l=0.186094u w=1.28u 
.ENDS senrq2

.SUBCKT seprq1 Q  CP D ENN SC SD SDN VDD VSS
MM56 IPS 5 13 VDD P l=0.18u w=0.52u 
MM42 VDD ENN 15 VDD P l=0.18u w=0.52u 
MM40 2 ENN VDD VDD P l=0.186783u w=1.15u 
MM38 VDD 16 2 VDD P l=0.186387u w=1.146u 
MM36 VDD SC 16 VDD P l=0.18u w=0.6u 
MM35 VDD SD 20 VDD P l=0.18u w=0.86u 
MM33 19 20 VDD VDD P l=0.18u w=0.98u 
MM32 24 16 30 VDD P l=0.18u w=0.52u 
MM34 VDD 19 30 VDD P l=0.18u w=0.52u 
MM31 VDD 16 22 VDD P l=0.18u w=0.64u 
MM60 VDD 2 21 VDD P l=0.18u w=0.52u 
MM59 VDD D 29 VDD P l=0.18u w=0.64u 
MM58 24 4 29 VDD P l=0.18u w=0.58u 
MM57 24 2 25 VDD P l=0.18u w=0.58u 
MM43 VDD 13 25 VDD P l=0.18u w=0.57u 
MM39 VDD 4 23 VDD P l=0.18u w=0.52u 
MM41 VDD 15 4 VDD P l=0.18u w=0.52u 
MM37 VDD 16 4 VDD P l=0.18u w=0.52u 
MM55 8 6 IPS VDD P l=0.18u w=0.52u 
MM54 6 CP VDD VDD P l=0.188434u w=1.245u 
MM53 VDD 6 5 VDD P l=0.18u w=1.26u 
MM51 24 5 IPM VDD P l=0.18u w=0.52u 
MM49 27 6 IPM VDD P l=0.18u w=0.61u 
MM52 VDD 8 27 VDD P l=0.18u w=0.61u 
MM50 8 IPM VDD VDD P l=0.18u w=1.19u 
MM48 8 SDN VDD VDD P l=0.187822u w=1.281u 
MM47 VDD IPS 12 VDD P l=0.18u w=0.63u 
MM46 Q 12 VDD VDD P l=0.18u w=1.5u 
MM45 VDD 12 13 VDD P l=0.18u w=0.59u 
MM44 13 SDN VDD VDD P l=0.18u w=0.59u 
MM19 IPS 5 8 VSS N l=0.18u w=0.44u 
MM18 33 IPM 8 VSS N l=0.18u w=0.82u 
MM9 2 ENN 32 VSS N l=0.18u w=0.49u 
MM12 VSS ENN 15 VSS N l=0.18u w=0.44u 
MM6 24 22 30 VSS N l=0.18u w=0.44u 
MM5 VSS 19 30 VSS N l=0.18u w=0.44u 
MM4 VSS 20 19 VSS N l=0.18u w=0.96u 
MM3 VSS 16 22 VSS N l=0.18u w=0.44u 
MM2 16 SC VSS VSS N l=0.18u w=0.65u 
MM1 20 SD VSS VSS N l=0.18u w=0.64u 
MM30 21 2 VSS VSS N l=0.18u w=0.44u 
MM29 24 21 25 VSS N l=0.18u w=0.44u 
MM28 24 23 29 VSS N l=0.18u w=0.44u 
MM27 29 D VSS VSS N l=0.18u w=0.44u 
MM11 23 4 VSS VSS N l=0.18u w=0.44u 
MM10 4 15 31 VSS N l=0.18u w=0.44u 
MM8 VSS 16 31 VSS N l=0.18u w=0.44u 
MM7 VSS 16 32 VSS N l=0.18u w=0.49u 
MM24 VSS 13 25 VSS N l=0.18u w=0.44u 
MM23 6 CP VSS VSS N l=0.186628u w=1.032u 
MM22 VSS 6 5 VSS N l=0.18u w=0.94u 
MM21 VSS 8 27 VSS N l=0.18u w=0.44u 
MM20 IPM 5 27 VSS N l=0.18u w=0.44u 
MM17 24 6 IPM VSS N l=0.18u w=0.44u 
MM13 VSS SDN 33 VSS N l=0.18u w=0.82u 
MM26 VSS IPS 12 VSS N l=0.18u w=0.52u 
MM25 VSS 12 Q VSS N l=0.18u w=1.08u 
MM16 13 6 IPS VSS N l=0.18u w=0.44u 
MM15 13 12 34 VSS N l=0.18u w=0.75u 
MM14 34 SDN VSS VSS N l=0.18u w=0.75u 
.ENDS seprq1

.SUBCKT seprq2 Q  CP D ENN SC SD SDN VDD VSS
MM58 IPS 5 13 VDD P l=0.18u w=0.52u 
MM43 VDD ENN 15 VDD P l=0.18u w=0.52u 
MM41 3 ENN VDD VDD P l=0.186783u w=1.15u 
MM39 VDD 16 3 VDD P l=0.186387u w=1.146u 
MM37 VDD SC 16 VDD P l=0.18u w=0.6u 
MM36 VDD SD 20 VDD P l=0.18u w=0.86u 
MM34 19 20 VDD VDD P l=0.18u w=0.98u 
MM33 24 16 30 VDD P l=0.18u w=0.52u 
MM35 VDD 19 30 VDD P l=0.18u w=0.52u 
MM32 VDD 16 22 VDD P l=0.18u w=0.64u 
MM62 VDD D 29 VDD P l=0.18u w=0.64u 
MM60 24 4 29 VDD P l=0.18u w=0.58u 
MM61 VDD 3 21 VDD P l=0.18u w=0.52u 
MM59 24 3 25 VDD P l=0.18u w=0.58u 
MM44 VDD 13 25 VDD P l=0.18u w=0.57u 
MM40 VDD 4 23 VDD P l=0.18u w=0.52u 
MM42 VDD 15 4 VDD P l=0.18u w=0.52u 
MM38 VDD 16 4 VDD P l=0.18u w=0.52u 
MM57 8 6 IPS VDD P l=0.18u w=0.52u 
MM56 6 CP VDD VDD P l=0.188434u w=1.245u 
MM55 VDD 6 5 VDD P l=0.18u w=1.26u 
MM53 24 5 IPM VDD P l=0.18u w=0.52u 
MM51 27 6 IPM VDD P l=0.18u w=0.61u 
MM54 VDD 8 27 VDD P l=0.18u w=0.61u 
MM52 8 IPM VDD VDD P l=0.18u w=1.19u 
MM50 8 SDN VDD VDD P l=0.187822u w=1.281u 
MM49 VDD IPS 12 VDD P l=0.18u w=0.63u 
MM48 VDD 12 Q VDD P l=0.18526u w=1.574u 
MM47 Q 12 VDD VDD P l=0.18u w=1.5u 
MM46 VDD 12 13 VDD P l=0.18u w=0.59u 
MM45 13 SDN VDD VDD P l=0.18u w=0.59u 
MM24 VSS 13 25 VSS N l=0.18u w=0.44u 
MM19 IPS 5 8 VSS N l=0.18u w=0.44u 
MM18 33 IPM 8 VSS N l=0.18u w=0.82u 
MM12 VSS ENN 15 VSS N l=0.18u w=0.44u 
MM9 3 ENN 32 VSS N l=0.18u w=0.49u 
MM6 VSS 16 22 VSS N l=0.18u w=0.44u 
MM5 16 SC VSS VSS N l=0.18u w=0.65u 
MM4 20 SD VSS VSS N l=0.18u w=0.64u 
MM3 24 22 30 VSS N l=0.18u w=0.44u 
MM2 VSS 19 30 VSS N l=0.18u w=0.44u 
MM1 VSS 20 19 VSS N l=0.18u w=0.96u 
MM31 24 21 25 VSS N l=0.18u w=0.44u 
MM30 24 23 29 VSS N l=0.18u w=0.44u 
MM29 29 D VSS VSS N l=0.18u w=0.44u 
MM28 21 3 VSS VSS N l=0.18u w=0.44u 
MM11 23 4 VSS VSS N l=0.18u w=0.44u 
MM10 4 15 31 VSS N l=0.18u w=0.44u 
MM8 VSS 16 31 VSS N l=0.18u w=0.44u 
MM7 VSS 16 32 VSS N l=0.18u w=0.49u 
MM23 6 CP VSS VSS N l=0.186628u w=1.032u 
MM22 VSS 6 5 VSS N l=0.18u w=0.94u 
MM21 VSS 8 27 VSS N l=0.18u w=0.44u 
MM20 IPM 5 27 VSS N l=0.18u w=0.44u 
MM17 24 6 IPM VSS N l=0.18u w=0.44u 
MM13 VSS SDN 33 VSS N l=0.18u w=0.82u 
MM27 VSS IPS 12 VSS N l=0.18u w=0.52u 
MM26 VSS 12 Q VSS N l=0.187175u w=1.154u 
MM25 VSS 12 Q VSS N l=0.18u w=1.08u 
MM16 13 6 IPS VSS N l=0.18u w=0.44u 
MM15 13 12 34 VSS N l=0.18u w=0.75u 
MM14 34 SDN VSS VSS N l=0.18u w=0.75u 
.ENDS seprq2

.SUBCKT srlab1 Q QN  RN SN VDD VSS
MM12 VDD 2 QN VDD P l=0.184785u w=1.63u 
MM11 5 2 VDD VDD P l=0.18671u w=1.234u 
MM9 5 RN VDD VDD P l=0.18u w=1.16u 
MM10 VDD SN 2 VDD P l=0.18u w=1.04u 
MM8 VDD 5 2 VDD P l=0.18u w=1.04u 
MM7 VDD 5 Q VDD P l=0.18u w=1.54u 
MM6 VSS 2 9 VSS N l=0.18u w=1.36u 
MM4 5 RN 9 VSS N l=0.18u w=1.36u 
MM3 10 5 2 VSS N l=0.18u w=1.36u 
MM5 10 SN VSS VSS N l=0.18u w=1.36u 
MM2 VSS 2 QN VSS N l=0.18u w=0.99u 
MM1 VSS 5 Q VSS N l=0.18u w=0.99u 
.ENDS srlab1

.SUBCKT srlab2 Q QN  RN SN VDD VSS
MM15 VDD 2 QN VDD P l=0.18427u w=1.602u 
MM14 VDD 2 QN VDD P l=0.18427u w=1.602u 
MM12 Q 3 VDD VDD P l=0.184324u w=1.582u 
MM11 Q 3 VDD VDD P l=0.184324u w=1.582u 
MM13 3 2 VDD VDD P l=0.18671u w=1.234u 
MM9 3 RN VDD VDD P l=0.18u w=1.16u 
MM10 VDD SN 2 VDD P l=0.18u w=1.04u 
MM8 VDD 3 2 VDD P l=0.18u w=1.04u 
MM7 QN 2 VSS VSS N l=0.185886u w=1.162u 
MM6 QN 2 VSS VSS N l=0.18u w=1.1u 
MM5 Q 3 VSS VSS N l=0.195401u w=1.87u 
MM4 VSS 2 9 VSS N l=0.18u w=1.36u 
MM2 3 RN 9 VSS N l=0.18u w=1.36u 
MM1 10 3 2 VSS N l=0.18u w=1.36u 
MM3 10 SN VSS VSS N l=0.18u w=1.36u 
.ENDS srlab2

.SUBCKT su01d0 CO S  A B CI VDD VSS
MM30 14 2 7 VDD P l=0.18u w=1.54u 
MM22 20 CI 7 VDD P l=0.18u w=1.2u 
MM29 VDD A 14 VDD P l=0.185695u w=1.454u 
MM18 VDD CI 14 VDD P l=0.18u w=1.22u 
MM28 19 A 2 VDD P l=0.18u w=1.38u 
MM19 13 CI 2 VDD P l=0.186047u w=1.29u 
MM26 14 4 VDD VDD P l=0.185697u w=1.622u 
MM27 20 A 18 VDD P l=0.18u w=1.2u 
MM25 VDD 4 18 VDD P l=0.18u w=1.2u 
MM23 19 4 VDD VDD P l=0.18u w=1.38u 
MM21 4 B VDD VDD P l=0.187374u w=1.188u 
MM20 13 A VDD VDD P l=0.186047u w=1.29u 
MM24 13 4 VDD VDD P l=0.18u w=1.22u 
MM16 S 7 VDD VDD P l=0.18u w=0.72u 
MM17 VDD 2 CO VDD P l=0.18u w=0.72u 
MM15 9 2 7 VSS N l=0.18u w=0.75u 
MM3 9 CI VSS VSS N l=0.18u w=0.58u 
MM12 15 A 17 VSS N l=0.18u w=0.75u 
MM11 VSS 4 15 VSS N l=0.18u w=0.75u 
MM14 16 A 2 VSS N l=0.18u w=1.22u 
MM9 16 4 VSS VSS N l=0.18u w=1.22u 
MM13 9 A VSS VSS N l=0.18u w=1.06u 
MM8 9 4 VSS VSS N l=0.187302u w=1.134u 
MM7 17 CI 7 VSS N l=0.18u w=0.75u 
MM6 VSS B 4 VSS N l=0.18u w=0.79u 
MM5 VSS A 12 VSS N l=0.186047u w=1.29u 
MM10 VSS 4 12 VSS N l=0.18u w=1.22u 
MM4 12 CI 2 VSS N l=0.186047u w=1.29u 
MM2 CO 2 VSS VSS N l=0.18u w=0.57u 
MM1 S 7 VSS VSS N l=0.18u w=0.57u 
.ENDS su01d0

.SUBCKT su01d1 CO S  A B CI VDD VSS
MM30 14 2 7 VDD P l=0.18u w=1.54u 
MM22 20 CI 7 VDD P l=0.18u w=1.2u 
MM29 VDD A 14 VDD P l=0.185695u w=1.454u 
MM18 VDD CI 14 VDD P l=0.18u w=1.22u 
MM28 19 A 2 VDD P l=0.18u w=1.38u 
MM19 13 CI 2 VDD P l=0.186047u w=1.29u 
MM26 14 4 VDD VDD P l=0.185697u w=1.622u 
MM27 20 A 18 VDD P l=0.18u w=1.2u 
MM25 VDD 4 18 VDD P l=0.18u w=1.2u 
MM23 19 4 VDD VDD P l=0.18u w=1.38u 
MM21 4 B VDD VDD P l=0.187374u w=1.188u 
MM20 13 A VDD VDD P l=0.186047u w=1.29u 
MM24 13 4 VDD VDD P l=0.18u w=1.22u 
MM17 VDD 2 CO VDD P l=0.18u w=1.55u 
MM16 VDD 7 S VDD P l=0.184815u w=1.62u 
MM15 9 2 7 VSS N l=0.18u w=0.75u 
MM3 9 CI VSS VSS N l=0.18u w=0.58u 
MM12 15 A 17 VSS N l=0.18u w=0.75u 
MM11 VSS 4 15 VSS N l=0.18u w=0.75u 
MM14 16 A 2 VSS N l=0.18u w=1.22u 
MM9 16 4 VSS VSS N l=0.18u w=1.22u 
MM13 9 A VSS VSS N l=0.18u w=1.06u 
MM8 9 4 VSS VSS N l=0.187302u w=1.134u 
MM7 17 CI 7 VSS N l=0.18u w=0.75u 
MM6 VSS B 4 VSS N l=0.18u w=0.79u 
MM5 VSS A 12 VSS N l=0.186047u w=1.29u 
MM10 VSS 4 12 VSS N l=0.18u w=1.22u 
MM4 12 CI 2 VSS N l=0.186047u w=1.29u 
MM2 CO 2 VSS VSS N l=0.187156u w=1.09u 
MM1 S 7 VSS VSS N l=0.18u w=1.12u 
.ENDS su01d1

.SUBCKT su01d2 CO S  A B CI VDD VSS
MM34 VDD A 13 VDD P l=0.185695u w=1.454u 
MM22 VDD CI 13 VDD P l=0.18u w=1.22u 
MM33 19 A 6 VDD P l=0.18u w=1.38u 
MM23 12 CI 6 VDD P l=0.186047u w=1.29u 
MM32 20 A 18 VDD P l=0.18u w=1.2u 
MM30 VDD 3 18 VDD P l=0.18u w=1.2u 
MM28 19 3 VDD VDD P l=0.18u w=1.38u 
MM27 3 B VDD VDD P l=0.187374u w=1.188u 
MM26 20 CI 7 VDD P l=0.18u w=1.2u 
MM25 12 A VDD VDD P l=0.186047u w=1.29u 
MM24 13 6 7 VDD P l=0.18u w=1.54u 
MM31 13 3 VDD VDD P l=0.185697u w=1.622u 
MM29 12 3 VDD VDD P l=0.18u w=1.22u 
MM21 VDD 6 CO VDD P l=0.185036u w=1.644u 
MM20 CO 6 VDD VDD P l=0.18u w=1.57u 
MM19 S 7 VDD VDD P l=0.185036u w=1.644u 
MM18 VDD 7 S VDD P l=0.18u w=1.57u 
MM15 15 A 17 VSS N l=0.18u w=0.75u 
MM14 VSS 3 15 VSS N l=0.18u w=0.75u 
MM17 16 A 6 VSS N l=0.18u w=1.22u 
MM12 16 3 VSS VSS N l=0.18u w=1.22u 
MM16 14 A VSS VSS N l=0.18u w=1.06u 
MM11 14 3 VSS VSS N l=0.187302u w=1.134u 
MM10 VSS B 3 VSS N l=0.18u w=0.95u 
MM9 17 CI 7 VSS N l=0.18u w=0.75u 
MM8 CO 6 VSS VSS N l=0.186935u w=1.194u 
MM7 CO 6 VSS VSS N l=0.18u w=1.12u 
MM6 S 7 VSS VSS N l=0.186935u w=1.194u 
MM5 VSS 7 S VSS N l=0.18u w=1.12u 
MM4 VSS A 11 VSS N l=0.186047u w=1.29u 
MM3 14 6 7 VSS N l=0.18u w=0.75u 
MM1 14 CI VSS VSS N l=0.18u w=0.58u 
MM13 VSS 3 11 VSS N l=0.18u w=1.22u 
MM2 11 CI 6 VSS N l=0.186047u w=1.29u 
.ENDS su01d2

.SUBCKT xn02d1 ZN  A1 A2 VDD VSS
MM13 4 A2 VDD VDD P l=0.18u w=0.55u 
MM12 5 A1 VDD VDD P l=0.18u w=0.63u 
MM11 11 A1 6 VDD P l=0.18u w=1.52u 
MM10 11 4 VDD VDD P l=0.18u w=1.52u 
MM14 VDD A2 12 VDD P l=0.184906u w=1.59u 
MM9 6 5 12 VDD P l=0.184906u w=1.59u 
MM8 VDD 6 ZN VDD P l=0.1852u w=1.5u 
MM7 6 A2 9 VSS N l=0.184465u w=1.532u 
MM2 6 5 10 VSS N l=0.18u w=1.03u 
MM6 4 A2 VSS VSS N l=0.18u w=0.48u 
MM5 9 A1 VSS VSS N l=0.184465u w=1.532u 
MM4 VSS A1 5 VSS N l=0.18u w=0.74u 
MM3 VSS 4 10 VSS N l=0.18u w=1.03u 
MM1 ZN 6 VSS VSS N l=0.18u w=1u 
.ENDS xn02d1

.SUBCKT xn02d2 ZN  A1 A2 VDD VSS
MM15 3 A2 VDD VDD P l=0.18u w=0.55u 
MM16 VDD A2 11 VDD P l=0.184906u w=1.59u 
MM13 6 4 11 VDD P l=0.184906u w=1.59u 
MM12 4 A1 VDD VDD P l=0.18u w=0.63u 
MM11 12 A1 6 VDD P l=0.18u w=1.52u 
MM14 12 3 VDD VDD P l=0.18u w=1.52u 
MM10 ZN 6 VDD VDD P l=0.185098u w=1.53u 
MM9 ZN 6 VDD VDD P l=0.18u w=1.46u 
MM8 6 A2 10 VSS N l=0.184465u w=1.532u 
MM5 6 4 9 VSS N l=0.18u w=1.03u 
MM7 3 A2 VSS VSS N l=0.18u w=0.48u 
MM6 VSS 3 9 VSS N l=0.18u w=1.03u 
MM4 10 A1 VSS VSS N l=0.184465u w=1.532u 
MM3 VSS A1 4 VSS N l=0.18u w=0.74u 
MM2 ZN 6 VSS VSS N l=0.186998u w=1.046u 
MM1 ZN 6 VSS VSS N l=0.18u w=0.98u 
.ENDS xn02d2

.SUBCKT xn02d4 ZN  A1 A2 VDD VSS
MM16 VDD A2 2 VDD P l=0.18u w=0.55u 
MM17 VDD A2 11 VDD P l=0.184906u w=1.59u 
MM15 6 4 11 VDD P l=0.185194u w=1.594u 
MM14 4 A1 VDD VDD P l=0.18u w=0.63u 
MM13 6 A1 12 VDD P l=0.18u w=1.52u 
MM18 VDD 2 12 VDD P l=0.18u w=1.52u 
MM12 ZN 6 VDD VDD P l=0.1839u w=2u 
MM11 ZN 6 VDD VDD P l=0.18u w=1.93u 
MM10 VDD 6 ZN VDD P l=0.183667u w=1.996u 
MM8 6 A2 10 VSS N l=0.185065u w=1.54u 
MM6 6 4 9 VSS N l=0.18u w=1.03u 
MM7 2 A2 VSS VSS N l=0.18u w=0.48u 
MM9 VSS 2 9 VSS N l=0.18u w=1.03u 
MM5 10 A1 VSS VSS N l=0.185065u w=1.54u 
MM4 VSS A1 4 VSS N l=0.18u w=0.74u 
MM3 ZN 6 VSS VSS N l=0.186161u w=1.344u 
MM2 VSS 6 ZN VSS N l=0.185821u w=1.34u 
MM1 ZN 6 VSS VSS N l=0.18u w=1.27u 
.ENDS xn02d4

.SUBCKT xr02d1 Z  A1 A2 VDD VSS
MM13 VDD A1 2 VDD P l=0.18u w=0.5u 
MM14 5 2 11 VDD P l=0.18u w=0.96u 
MM12 12 A1 5 VDD P l=0.18u w=0.96u 
MM11 11 4 VDD VDD P l=0.18u w=0.96u 
MM10 Z 5 VDD VDD P l=0.186152u w=1.502u 
MM9 VDD A2 4 VDD P l=0.18u w=0.48u 
MM8 VDD A2 12 VDD P l=0.18u w=0.96u 
MM7 9 2 5 VSS N l=0.18u w=0.59u 
MM1 VSS A2 9 VSS N l=0.18u w=0.52u 
MM5 10 A1 5 VSS N l=0.18u w=0.67u 
MM6 VSS A1 2 VSS N l=0.18u w=0.48u 
MM4 VSS 4 10 VSS N l=0.18u w=0.67u 
MM3 VSS 5 Z VSS N l=0.187349u w=0.996u 
MM2 VSS A2 4 VSS N l=0.18u w=0.48u 
.ENDS xr02d1

.SUBCKT xr02d2 Z  A1 A2 VDD VSS
MM15 VDD A1 2 VDD P l=0.18u w=0.5u 
MM16 5 2 11 VDD P l=0.18u w=0.96u 
MM14 12 A1 5 VDD P l=0.18u w=0.96u 
MM13 11 4 VDD VDD P l=0.18u w=0.96u 
MM12 Z 5 VDD VDD P l=0.186152u w=1.502u 
MM11 Z 5 VDD VDD P l=0.186152u w=1.502u 
MM10 VDD A2 4 VDD P l=0.18u w=0.48u 
MM9 VDD A2 12 VDD P l=0.18u w=0.96u 
MM8 9 2 5 VSS N l=0.18u w=0.59u 
MM1 VSS A2 9 VSS N l=0.18u w=0.52u 
MM6 5 A1 10 VSS N l=0.18u w=0.67u 
MM7 VSS A1 2 VSS N l=0.18u w=0.48u 
MM5 VSS 4 10 VSS N l=0.18u w=0.67u 
MM4 VSS 5 Z VSS N l=0.187349u w=0.996u 
MM3 VSS 5 Z VSS N l=0.187349u w=0.996u 
MM2 VSS A2 4 VSS N l=0.18u w=0.48u 
.ENDS xr02d2

.SUBCKT xr02d4 Z  A1 A2 VDD VSS
MM18 VDD A1 5 VDD P l=0.18u w=0.5u 
MM15 VDD 4 Z VDD P l=0.189022u w=2.168u 
MM14 VDD 4 Z VDD P l=0.185911u w=2.101u 
MM13 Z 4 VDD VDD P l=0.18u w=1.59u 
MM16 11 3 VDD VDD P l=0.18u w=0.96u 
MM12 4 5 11 VDD P l=0.18u w=0.96u 
MM17 12 A1 4 VDD P l=0.18u w=0.96u 
MM11 VDD A2 3 VDD P l=0.18u w=0.48u 
MM10 VDD A2 12 VDD P l=0.18u w=0.96u 
MM9 VSS A1 5 VSS N l=0.18u w=0.48u 
MM8 4 A1 9 VSS N l=0.18u w=0.67u 
MM3 10 5 4 VSS N l=0.18u w=0.59u 
MM7 VSS 3 9 VSS N l=0.18u w=0.67u 
MM6 VSS 4 Z VSS N l=0.189333u w=1.125u 
MM5 VSS 4 Z VSS N l=0.186679u w=1.096u 
MM4 VSS 4 Z VSS N l=0.184643u w=1.68u 
MM1 VSS A2 10 VSS N l=0.18u w=0.52u 
MM2 VSS A2 3 VSS N l=0.18u w=0.48u 
.ENDS xr02d4

.SUBCKT xr03d1 Z  A1 A2 A3 VDD VSS
MM22 10 2 VDD VDD P l=0.18u w=0.64u 
MM21 VDD A3 4 VDD P l=0.186564u w=1.042u 
MM19 2 A2 4 VDD P l=0.18u w=0.98u 
MM18 6 A2 VDD VDD P l=0.18u w=0.98u 
MM20 14 4 VDD VDD P l=0.18u w=0.98u 
MM17 14 6 2 VDD P l=0.18u w=0.98u 
MM15 VDD 7 Z VDD P l=0.184554u w=1.502u 
MM16 13 2 7 VDD P l=0.18u w=1.54u 
MM14 VDD 8 13 VDD P l=0.18427u w=1.602u 
MM13 VDD A1 8 VDD P l=0.184845u w=1.61u 
MM12 7 10 8 VDD P l=0.18u w=1.54u 
MM11 VSS 2 10 VSS N l=0.18u w=0.54u 
MM8 VSS A2 6 VSS N l=0.18u w=0.75u 
MM9 VSS 4 14 VSS N l=0.18u w=0.75u 
MM7 14 A2 2 VSS N l=0.18u w=0.75u 
MM6 4 6 2 VSS N l=0.18u w=0.75u 
MM10 4 A3 VSS VSS N l=0.18u w=0.75u 
MM5 8 2 7 VSS N l=0.18u w=1.23u 
MM4 8 A1 VSS VSS N l=0.18u w=0.72u 
MM3 VSS 7 Z VSS N l=0.18u w=1u 
MM2 VSS 8 13 VSS N l=0.18635u w=1.304u 
MM1 13 10 7 VSS N l=0.18u w=1.23u 
.ENDS xr03d1

.SUBCKT xr03d2 Z  A1 A2 A3 VDD VSS
MM24 7 2 VDD VDD P l=0.18u w=0.64u 
MM23 VDD A3 4 VDD P l=0.186564u w=1.042u 
MM21 2 A2 4 VDD P l=0.18u w=0.98u 
MM20 6 A2 VDD VDD P l=0.18u w=0.98u 
MM22 14 4 VDD VDD P l=0.18u w=0.98u 
MM19 14 6 2 VDD P l=0.18u w=0.98u 
MM18 8 7 9 VDD P l=0.18u w=1.54u 
MM17 13 2 8 VDD P l=0.18u w=1.54u 
MM16 VDD 8 Z VDD P l=0.184554u w=1.502u 
MM15 VDD 8 Z VDD P l=0.184554u w=1.502u 
MM14 VDD 9 13 VDD P l=0.18427u w=1.602u 
MM13 VDD A1 9 VDD P l=0.184845u w=1.61u 
MM11 9 2 8 VSS N l=0.18u w=1.23u 
MM10 9 A1 VSS VSS N l=0.18u w=0.72u 
MM12 13 7 8 VSS N l=0.18u w=1.23u 
MM9 VSS 8 Z VSS N l=0.186826u w=1.002u 
MM8 VSS 8 Z VSS N l=0.18u w=1u 
MM7 VSS 9 13 VSS N l=0.18635u w=1.304u 
MM6 VSS 2 7 VSS N l=0.18u w=0.54u 
MM3 VSS A2 6 VSS N l=0.18u w=0.75u 
MM4 VSS 4 14 VSS N l=0.18u w=0.75u 
MM2 14 A2 2 VSS N l=0.18u w=0.75u 
MM1 4 6 2 VSS N l=0.18u w=0.75u 
MM5 4 A3 VSS VSS N l=0.18u w=0.75u 
.ENDS xr03d2

.SUBCKT xr03d4 Z  A1 A2 A3 VDD VSS
MM26 VDD A1 5 VDD P l=0.184845u w=1.61u 
MM25 6 3 5 VDD P l=0.18u w=1.54u 
MM24 13 4 6 VDD P l=0.18u w=1.54u 
MM23 VDD 5 13 VDD P l=0.18427u w=1.602u 
MM22 Z 6 VDD VDD P l=0.187066u w=2.072u 
MM21 Z 6 VDD VDD P l=0.186277u w=2.055u 
MM20 VDD 6 Z VDD P l=0.18688u w=1.875u 
MM19 3 4 VDD VDD P l=0.18u w=0.64u 
MM18 VDD A3 8 VDD P l=0.186564u w=1.042u 
MM16 4 A2 8 VDD P l=0.18u w=0.98u 
MM15 10 A2 VDD VDD P l=0.18u w=0.98u 
MM17 14 8 VDD VDD P l=0.18u w=0.98u 
MM14 14 10 4 VDD P l=0.18u w=0.98u 
MM12 5 4 6 VSS N l=0.18u w=1.23u 
MM11 5 A1 VSS VSS N l=0.18u w=0.72u 
MM13 13 3 6 VSS N l=0.18u w=1.23u 
MM10 VSS 5 13 VSS N l=0.18635u w=1.304u 
MM8 Z 6 VSS VSS N l=0.185097u w=1.342u 
MM9 VSS 6 Z VSS N l=0.185022u w=1.362u 
MM7 VSS 6 Z VSS N l=0.18u w=1.3u 
MM6 VSS 4 3 VSS N l=0.18u w=0.54u 
MM3 VSS A2 10 VSS N l=0.18u w=0.75u 
MM4 VSS 8 14 VSS N l=0.18u w=0.75u 
MM2 14 A2 4 VSS N l=0.18u w=0.75u 
MM1 8 10 4 VSS N l=0.18u w=0.75u 
MM5 8 A3 VSS VSS N l=0.18u w=0.75u 
.ENDS xr03d4

.SUBCKT ad01d4 CO S  A B CI VDD VSS
M1      U50_drain CI      U50_source VSS     N   L=0.18U  W=0.55U  
M2      U48_drain B       VSS     VSS     N   L=0.18U  W=0.65U  
M3      U68_in  CI      u12_source VSS     N   L=0.18U  W=0.65U  
M4      u12_source B       VSS     VSS     N   L=0.18U  W=0.69U  
M5      u12_source A       VSS     VSS     N   L=0.18U  W=0.69U  
M6      U68_in  A       U48_drain VSS     N   L=0.18U  W=0.65U  
M7      U50_drain U68_in  U53_source VSS     N   L=0.18U  W=0.55U  
M8      U53_source B       VSS     VSS     N   L=0.18U  W=0.55U  
M9      U53_source A       VSS     VSS     N   L=0.18U  W=0.55U  
M10     U53_source CI      VSS     VSS     N   L=0.18U  W=0.55U  
M11     U50_source A       U51_source VSS     N   L=0.18U  W=0.55U  
M12     U51_source B       VSS     VSS     N   L=0.18U  W=0.55U  
M13     S       U50_drain VSS     VSS     N   L=0.18U  W=2.94U  
M14     S       U50_drain VDD     VDD     P   L=0.182U  W=8.58U  
M15     CO      U68_in  VSS     VSS     N   L=0.18U  W=2.94U  
M16     CO      U68_in  VDD     VDD     P   L=0.184U  W=8.38U  
M17     U50_drain CI      U38_source VDD     P   L=0.185U  W=1.43U  
M18     u4_drain A       VDD     VDD     P   L=0.184U  W=1.77U  
M19     U68_in  CI      u4_drain VDD     P   L=0.185U  W=1.65U  
M20     u4_drain B       VDD     VDD     P   L=0.18U  W=1.77U  
M21     U41_drain B       VDD     VDD     P   L=0.185U  W=1.65U  
M22     U68_in  A       U41_drain VDD     P   L=0.185U  W=1.65U  
M23     U33_drain CI      VDD     VDD     P   L=0.18U  W=1.43U  
M24     U33_drain B       VDD     VDD     P   L=0.18U  W=1.41U  
M25     U50_drain U68_in  U33_drain VDD     P   L=0.185U  W=1.38U  
M26     U33_drain A       VDD     VDD     P   L=0.185U  W=1.43U  
M27     U38_source A       U37_source VDD     P   L=0.185U  W=1.43U  
M28     U37_source B       VDD     VDD     P   L=0.185U  W=1.43U  

.ENDS ad01d4

.SUBCKT adp1d4 CO P S  A B CI VDD VSS
M1      U63_drain U63_gate U63_source VSS     N   L=0.18U   W=0.55U
M2      U29_drain A       U29_source VSS     N   L=0.18U    W=0.55U
M3      U63_source B       VSS     VSS     N   L=0.18U     W=0.55U
M4      U29_source B       VSS     VSS     N   L=0.18U    W=0.55U
M5      U29_drain U30_gate U31_source VSS     N   L=0.18U    W=0.55U
M6      U31_source CI      VSS     VSS     N   L=0.18U     W=0.55U
M7      U56_drain A       VSS     VSS     N   L=0.18U    W=0.55U
M8      U63_drain U61_gate U56_drain VSS     N   L=0.18U    W=0.55U
M9      u13_drain CI      VSS     VSS     N   L=0.18U      W=0.61U
M10     u5_source U63_drain u13_drain VSS     N   L=0.18U    W=0.61U
M11     u11_drain U54_out VSS     VSS     N   L=0.18U    W=0.61U
M12     u5_source U30_gate u11_drain VSS     N   L=0.18U      W=0.61U
M13     U30_drain U30_gate U29_drain VDD     P   L=0.185U     W=1.51U
M14     VDD     U61_gate U61_source VDD     P   L=0.18U     W=0.89U
M15     U61_source U63_gate U63_drain VDD     P   L=0.18U      W=0.89U
M16     VDD     B       U30_drain VDD     P   L=0.18U     W=1.51U
M17     U29_drain CI      U30_drain VDD     P   L=0.18U     W=1.51U
M18     U30_drain A       VDD     VDD     P   L=0.18U    W=1.51U
M19     U63_drain A       U64_source VDD     P   L=0.18U      W=1.16U
M20     U64_source B       VDD     VDD     P   L=0.18U      W=1.16U
M21     u2_drain CI      VDD     VDD     P   L=0.18U      W=1.56U
M22     u5_drain U63_drain u5_source VDD     P   L=0.187U    W=1.56U
M23     VDD     U54_out u5_drain VDD     P   L=0.187U     W=1.56U
M24     u5_source U30_gate u2_drain VDD     P   L=0.18U      W=1.56U
M25     U30_gate U63_drain VSS     VSS     N   L=0.18U     W=0.61U
M26     U30_gate U63_drain VDD     VDD     P   L=0.187U     W=1.56U
M27     U63_gate A       VSS     VSS     N   L=0.18U     W=0.55U
M28     U63_gate A       VDD     VDD     P   L=0.185U    W=1.51U
M29     U54_out CI      VSS     VSS     N   L=0.18U      W=0.58U
M30     U54_out CI      VDD     VDD     P   L=0.18U      W=1.56U
M31     U61_gate B       VSS     VSS     N   L=0.18U     W=0.55U
M32     U61_gate B       VDD     VDD     P   L=0.18U     W=1.52U
M33     CO      U29_drain VSS     VSS     N   L=0.184U    W=2.94U
M34     CO      U29_drain VDD     VDD     P   L=0.182U      W=8.56U
M35     P       U63_drain VSS     VSS     N   L=0.18U    W=3.07U
M36     P       U63_drain VDD     VDD     P   L=0.182U    W=8.28U
M37     S       u5_source VSS     VSS     N   L=0.182U     W=2.94U
M38     S       u5_source VDD     VDD     P   L=0.18U      W=8.64U

.ENDS adp1d4

.SUBCKT ah01d4 CO S  A B VDD VSS
M1      CO      U1_in   VSS     VSS       N   L=0.185U      W=2.91U
M2      CO      U1_in   VDD     VDD       P   L=0.185U      W=8.46U
M3      S       U5_in   VSS     VSS       N   L=0.183U      W=2.91U
M4      S       U5_in   VDD     VDD       P   L=0.184U      W=8.28U
M5      U1_in   A       VDD     VDD       P   L=0.184U      W=1.80U
M6      U1_in   B       VDD     VDD       P   L=0.184U      W=1.80U
M7      U5_in   A       U9_source VDD     P   L=0.18U       W=1.20U
M8      U9_source B       VDD     VDD     P   L=0.18U       W=1.20U
M9      U5_in   U1_in   VDD     VDD       P   L=0.18U       W=1.20U
M10     U75_drain B       VSS     VSS     N   L=0.18U       W=0.72U
M11     U1_in   A       U75_drain VSS     N   L=0.18U       W=0.72U
M12     U5_in   U1_in   U12_source VSS    N   L=0.18U       W=0.73U
M13     U12_source B       VSS     VSS    N   L=0.18U       W=0.39U
M14     U12_source A       VSS     VSS    N   L=0.18U       W=0.39U

.ENDS ah01d4

.SUBCKT an02d7 Z  A1 A2 VDD VSS
M1      U3_drain A2      VDD     VDD     P   L=0.184U  W=1.86U   
+  PD=.820U
M2      U3_drain A1      VDD     VDD     P   L=0.184U  W=1.86U   
+  PD=.820U
M3      Z       U3_drain VDD     VDD     P   L=0.185167U  W=14.37U   
+  PD=1.505U
M4      u2_drain A2      VSS     VSS     N   L=0.18U  W=1.01U   
+  PD=.700U
M5      U3_drain A1      u2_drain VSS     N   L=0.188U  W=1.01U   
+  PS=.700U PD=.700U
M6      Z       U3_drain VSS     VSS     N   L=0.18U  W=5.05U   
+  PD=1.382U

.ENDS an02d7

.SUBCKT an02da Z  A1 A2 VDD VSS
M1      U3_drain A2      VDD     VDD     P   L=0.18U       W=1.7U
+  PD=.820U
M2      U3_drain A1      VDD     VDD     P   L=0.185U      W=1.7U
+  PD=.820U
M3      Z       U3_drain VDD     VDD     P   L=0.18275U      W=20.22U
+  PD=1.505U
M4      u2_drain A2      VSS     VSS     N   L=0.18U       W=0.95U
+  PD=.700U
M5      U3_drain A1      u2_drain VSS     N   L=0.18U       W=0.95U
+  PS=.700U PD=.700U
M6      Z       U3_drain VSS     VSS     N   L=0.185U       W=7.42U
+  PD=1.382U

.ENDS an02da

.SUBCKT an03d7 Z  A1 A2 A3 VDD VSS
M1      U5_drain A3      VDD     VDD     P   L=0.185U  W=1.7U     
+  PD=.863U
M2      U5_drain A2      VDD     VDD     P   L=0.18U  W=1.7U     
+  PD=.863U
M3      U5_drain A1      VDD     VDD     P   L=0.184U  W=1.7U     
+  PD=.863U
M4      Z       U5_drain VDD     VDD     P   L=0.183U  W=14.51U     
+  PD=1.561U
M5      Z       U5_drain VSS     VSS     N   L=0.18U  W=4.98U     
+  PD=1.174U
M6      U5_drain A1      U4_source VSS     N   L=0.18U  W=0.95U     
+  PS=.890U PD=.890U
M7      U4_source A2      u2_source VSS     N   L=0.18U  W=0.95U     
+  PS=.890U PD=.890U
M8      u2_source A3      VSS     VSS     N   L=0.18U  W=0.95U     
+  PD=.890U

.ENDS an03d7

.SUBCKT an03da Z  A1 A2 A3 VDD VSS
M1      U5_drain A3      VDD     VDD     P   L=0.184U  W=1.7U     
+  PD=.863U
M2      U5_drain A2      VDD     VDD     P   L=0.184U  W=1.7U     
+  PD=.863U
M3      U5_drain A1      VDD     VDD     P   L=0.185U  W=1.7U     
+  PD=.863U
M4      Z       U5_drain VDD     VDD     P   L=0.183125U  W=19.99U     
+  PD=1.561U
M5      Z       U5_drain VSS     VSS     N   L=0.18U  W=7.53U     
+  PD=1.174U
M6      U5_drain A1      U4_source VSS     N   L=0.18U  W=0.87U    
+  PS=.890U PD=.890U
M7      U4_source A2      u2_source VSS     N   L=0.18U  W=0.87U     
+  PS=.890U PD=.890U
M8      u2_source A3      VSS     VSS     N   L=0.18U  W=0.87U     
+  PD=.890U

.ENDS an03da

.SUBCKT an04d7 Z  A1 A2 A3 A4 VDD VSS
M1      VDD     A4      U7_source VDD     P   L=0.185U  W=1.7U
+  PS=.875U
M2      VDD     A3      U7_source VDD     P   L=0.18U  W=1.7U
+  PS=.875U
M3      VDD     A2      U7_source VDD     P   L=0.185U  W=1.7U
+  PS=.875U
M4      VDD     A1      U7_source VDD     P   L=0.185U  W=1.7U
+  PS=.875U
M5      VDD     U7_source Z       VDD     P   L=0.182833U  W=14.51U
+  PS=1.496U
M6      Z       U7_source VSS     VSS     N   L=0.18U  W=5.05U
+  PD=1.054U
M7      u2_drain A2      u2_source VSS     N   L=0.18U  W=0.95U
+  PS=.900U PD=.900U
M8      u2_source A3      U6_source VSS     N   L=0.18U  W=0.95U
+  PS=.900U PD=.900U
M9      U6_source A4      VSS     VSS     N   L=0.18U  W=0.95U
+  PD=.900U
M10     U7_source A1      u2_drain VSS     N   L=0.18U  W=0.95U
+  PS=.900U PD=.900U

.ENDS an04d7

.SUBCKT an04da Z  A1 A2 A3 A4 VDD VSS
M1      VDD     A4      U7_source VDD     P   L=0.185U  W=1.7U
+  PS=.875U
M2      VDD     A3      U7_source VDD     P   L=0.18U  W=1.7U
+  PS=.875U
M3      VDD     A2      U7_source VDD     P   L=0.185U  W=1.7U
+  PS=.875U
M4      VDD     A1      U7_source VDD     P   L=0.185U  W=1.7U
+  PS=.875U
M5      VDD     U7_source Z       VDD     P   L=0.184U  W=17.83U
+  PS=1.496U
M6      Z       U7_source VSS     VSS     N   L=0.18U  W=7.42U
+  PD=1.054U
M7      u2_drain A2      u2_source VSS     N   L=0.18U  W=0.87U
+  PS=.900U PD=.900U
M8      u2_source A3      U6_source VSS     N   L=0.18U  W=0.87U
+  PS=.900U PD=.900U
M9      U6_source A4      VSS     VSS     N   L=0.18U  W=0.87U
+  PD=.900U
M10     U7_source A1      u2_drain VSS     N   L=0.18U  W=0.87U
+  PS=.900U PD=.900U

.ENDS an04da

.SUBCKT bufbd2 Z  I VDD VSS
M1      Z       U2_gate VDD     VDD     P   L=0.184U      W=4.1U
M2      U2_gate I       VDD     VDD     P   L=0.18U      W=2.19U
M3      Z       U2_gate VSS     VSS     N   L=0.18U      W=1.45U
M4      U2_gate I       VSS     VSS     N   L=0.18U      W=0.62U

.ENDS bufbd2

.SUBCKT bufbd4 Z  I VDD VSS
M1      Z       U2_gate VDD     VDD     P   L=0.182667U  W=7.27U  
M2      U2_gate I       VDD     VDD     P   L=0.1835U    W=2.26U  
M3      Z       U2_gate VSS     VSS     N   L=0.18U      W=2.91U  
M4      U2_gate I       VSS     VSS     N   L=0.18U      W=0.69U  

.ENDS bufbd4

.SUBCKT bufbdf Z  I VDD VSS
M1      Z       U2_gate VDD     VDD     P   L=0.183U  W=30.43U  
M2      U2_gate I       VDD     VDD     P   L=0.183U  W=5.03U  
M3      Z       U2_gate VSS     VSS     N   L=0.18U  W=10.76U  
M4      U2_gate I       VSS     VSS     N   L=0.18U  W=1.41U  

.ENDS bufbdf

.SUBCKT bufbdk Z  I VDD VSS
M1      Z       U2_gate VDD     VDD     P   L=0.182812U    W=40.68U
M2      U2_gate I       VDD     VDD     P   L=0.183333U     W=5.03U
M3      Z       U2_gate VSS     VSS     N   L=0.18U     W=14.41U
M4      U2_gate I       VSS     VSS     N   L=0.18U      W=1.41U

.ENDS bufbdk

.SUBCKT buffd2 Z  I VDD VSS
M1      Z       U39_gate VSS     VSS     N   L=0.18U      W=1.45U
M2      U39_gate I       VSS     VSS     N   L=0.18U      W=0.62U
M3      Z       U39_gate VDD     VDD     P   L=0.186U     W=4.16U
M4      U39_gate I       VDD     VDD     P   L=0.184U      W=1.76U

.ENDS buffd2

.SUBCKT buffd4 Z  I VDD VSS
M1      Z       U39_gate VSS     VSS     N   L=0.18U  W=2.91U  
M2      U39_gate I       VSS     VSS     N   L=0.18U  W=0.93U  
M3      Z       U39_gate VDD     VDD     P   L=0.1835U  W=8.49U  
M4      U39_gate I       VDD     VDD     P   L=0.1835U  W=2.26U  

.ENDS buffd4

.SUBCKT cg01d4 CO  A B CI VDD VSS
M1      CO      U68_in  VSS     VSS     N   L=0.18U  W=2.95U  
M2      CO      U68_in  VDD     VDD     P   L=0.184U  W=8.38U  
M3      U68_in  A       U42_source VDD     P   L=0.18U  W=1.87U  
M4      U68_in  CI      U32_source VDD     P   L=0.18U  W=1.87U  
M5      U32_source B       VDD     VDD     P   L=0.18U  W=1.87U  
M6      U32_source A       VDD     VDD     P   L=0.18U  W=1.87U  
M7      U42_source B       VDD     VDD     P   L=0.18U  W=1.87U  
M8      U68_in  A       U49_source VSS     N   L=0.18U  W=0.65U  
M9      U49_source B       VSS     VSS     N   L=0.18U  W=0.65U  
M10     U46_drain A       VSS     VSS     N   L=0.18U  W=0.65U  
M11     U46_drain B       VSS     VSS     N   L=0.18U  W=0.65U  
M12     U68_in  CI      U46_drain VSS     N   L=0.18U  W=0.65U  

.ENDS cg01d4

.SUBCKT decfq4 Q  CDN CPN D ENN VDD VSS
M1      U32_u7_drain CDN     VSS          VSS     N   L=0.18U   W=0.89U   
+  PD=.550U
M2      U32_out      U32_in1 U32_u7_drain VSS     N   L=0.18U   W=0.89U   
+  PS=.550U PD=.550U 
M3      U32_out      U32_in1 VDD          VDD     P   L=0.18U   W=1.29U   PD=.548U
M4      VDD          CDN     U32_out      VDD     P   L=0.186U  W=1.29U   PS=.548U
M5      U31_u7_drain CDN     VSS          VSS     N   L=0.18U   W=0.9U   
+  PD=.960U
M6      U23_in       u8_S    U31_u7_drain VSS     N   L=0.18U   W=0.9U   
+  PS=.960U PD=.960U
M7      U23_in       u8_S    VDD          VDD     P   L=0.184U  W=1.67U   PD=.960U
M8      VDD          CDN     U23_in       VDD     P   L=0.184U  W=1.67U   PS=.960U
M9      u8_S         u8_GB   U32_in1      VDD     P   L=0.186U  W=1.11U  
M10     u8_S         u8_G    U32_in1      VSS     N   L=0.18U   W=0.48U  
M11     U32_out      u8_GB   U22_in       VDD     P   L=0.186U  W=1.11U   PD=.548U
M12     U32_out      u8_G    U22_in       VSS     N   L=0.18U   W=0.44U   PD=.550U
M13     U22_in       u8_G    U15_D        VDD     P   L=0.18U   W=1.11U  
M14     U22_in       u8_GB   U15_D        VSS     N   L=0.18U   W=0.44U  
M15     U15_D        U30_out U28_D        VDD     P   L=0.18U   W=1.45U  
M16     U15_D        U30_in  U28_D        VSS     N   L=0.18U   W=0.62U  
M17     U15_D        U30_in  U27_D        VDD     P   L=0.18U   W=1.45U  
M18     U15_D        U30_out U27_D        VSS     N   L=0.18U   W=0.62U  
M19     U23_out      u8_G    u8_S         VDD     P   L=0.18U   W=1.11U  
M20     U23_out      u8_GB   u8_S         VSS     N   L=0.18U   W=0.48U  
M21     U32_in1      U22_in  VSS          VSS     N   L=0.18U   W=0.84U  
M22     U32_in1      U22_in  VDD          VDD     P   L=0.18U   W=1.66U  
M23     u8_G         CPN     VSS          VSS     N   L=0.18U   W=0.69U  
M24     u8_G         CPN     VDD          VDD     P   L=0.183U  W=2.01U  
M25     u8_GB        u8_G    VSS          VSS     N   L=0.18U   W=0.44U  
M26     u8_GB        u8_G    VDD          VDD     P   L=0.18U   W=1.25U  
M27     U30_out      U30_in  VSS          VSS     N   L=0.18U   W=0.62U  
M28     U30_out      U30_in  VDD          VDD     P   L=0.18U   W=1.55U  
M29     U30_in       ENN     VSS          VSS     N   L=0.18U   W=0.62U  
M30     U30_in       ENN     VDD          VDD     P   L=0.185U  W=1.55U  
M31     U28_D        D       VSS          VSS     N   L=0.18U   W=0.62U  
M32     U28_D        D       VDD          VDD     P   L=0.186U  W=1.55U  
M33     U23_out      U23_in  VSS          VSS     N   L=0.18U   W=0.72U  
M34     U23_out      U23_in  VDD          VDD     P   L=0.185U  W=1.48U  
M35     U27_D        U23_out VSS          VSS     N   L=0.18U  W=0.62U  
M36     U27_D        U23_out VDD          VDD     P   L=0.185U  W=1.45U  
M37     Q            U23_in  VSS          VSS     N   L=0.18U  W=2.91U  
M38     Q            U23_in  VDD          VDD     P   L=0.18U  W=8.28U  

.ENDS decfq4

.SUBCKT decrq4 Q  CDN CP D ENN VDD VSS
M1      U32_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.89U   
+  PD=.600U
M2      U32_out U32_in1 U32_u7_drain VSS     N   L=0.18U  W=0.89U   
+  PS=.600U PD=.600U
M3      U32_out U32_in1 VDD     VDD     P   L=0.18U  W=1.29U   PD=.600U
M4      VDD     CDN     U32_out VDD     P   L=0.186U  W=1.29U   PS=.600U
M5      U31_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.93U   
+  PD=1.000U
M6      U31_out u8_S    U31_u7_drain VSS     N   L=0.18U  W=0.93U   
+  PS=1.000U PD=1.000U
M7      U31_out u8_S    VDD     VDD     P   L=0.184U  W=1.66U   
+  PD=1.045U
M8      VDD     CDN     U31_out VDD     P   L=0.184U  W=1.66U   
+  PS=1.045U
M9      u8_S    u8_GB   U32_in1 VDD     P   L=0.186U  W=1.11U  
M10     u8_S    u8_G    U32_in1 VSS     N   L=0.18U  W=0.48U  
M11     U32_out u8_GB   U22_in  VDD     P   L=0.186U  W=1.11U   PD=.600U
M12     U32_out u8_G    U22_in  VSS     N   L=0.18U  W=0.48U   PD=.600U
M13     U28_S   U30_out U28_D   VDD     P   L=0.18U  W=1.45U  
M14     U28_S   U30_in  U28_D   VSS     N   L=0.18U  W=0.62U  
M15     U28_S   u8_G    U22_in  VDD     P   L=0.18U  W=1.11U  
M16     U28_S   u8_GB   U22_in  VSS     N   L=0.18U  W=0.48U  
M17     U28_S   U30_in  U27_D   VDD     P   L=0.18U  W=1.45U  
M18     U28_S   U30_out U27_D   VSS     N   L=0.18U  W=0.62U  
M19     U23_out u8_G    u8_S    VDD     P   L=0.18U  W=1.11U  
M20     U23_out u8_GB   u8_S    VSS     N   L=0.18U  W=0.48U  
M21     U32_in1 U22_in  VSS     VSS     N   L=0.18U  W=0.79U  
M22     U32_in1 U22_in  VDD     VDD     P   L=0.18U  W=1.66U  
M23     u8_G    u8_GB   VSS     VSS     N   L=0.18U  W=0.47U 
M24     u8_G    u8_GB   VDD     VDD     P   L=0.18U  W=1.38U  
M25     u8_GB   CP      VSS     VSS     N   L=0.18U  W=0.69U  
M26     u8_GB   CP      VDD     VDD     P   L=0.183U  W=1.88U  
M27     U30_out U30_in  VSS     VSS     N   L=0.18U  W=0.62U  
M28     U30_out U30_in  VDD     VDD     P   L=0.18U  W=1.55U  
M29     U30_in  ENN     VSS     VSS     N   L=0.18U  W=0.62U  
M30     U30_in  ENN     VDD     VDD     P   L=0.185U  W=1.55U  
M31     U28_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M32     U28_D   D       VDD     VDD     P   L=0.186U  W=1.55U  
M33     U23_out U31_out VSS     VSS     N   L=0.18U  W=0.72U  
M34     U23_out U31_out VDD     VDD     P   L=0.185U  W=1.48U  
M35     Q       U31_out VSS     VSS     N   L=0.18U  W=2.94U  
M36     Q       U31_out VDD     VDD     P   L=0.183U  W=8.2U  
M37     U27_D   U23_out VSS     VSS     N   L=0.18U  W=0.62U  
M38     U27_D   U23_out VDD     VDD     P   L=0.184U  W=1.52U  

.ENDS decrq4

.SUBCKT denrq4 Q  CP D ENN VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.187U  W=1.11U  
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U  W=0.48U  
M3      U24_out u8_GB   U22_in  VDD     P   L=0.18U  W=1.11U  
M4      U24_out u8_G    U22_in  VSS     N   L=0.18U  W=0.53U  
M5      U28_S   U28_GB  U28_D   VDD     P   L=0.18U  W=1.45U  
M6      U28_S   U28_G   U28_D   VSS     N   L=0.18U  W=0.62U  
M7      U28_S   U28_G   U27_D   VDD     P   L=0.185U  W=1.45U  
M8      U28_S   U28_GB  U27_D   VSS     N   L=0.18U  W=0.62U  
M9      U28_S   u8_G    U22_in  VDD     P   L=0.187U  W=1.11U  
M10     U28_S   u8_GB   U22_in  VSS     N   L=0.18U  W=0.53U  
M11     u9_S    u8_G    u8_S    VDD     P   L=0.187U  W=1.11U  
M12     u9_S    u8_GB   u8_S    VSS     N   L=0.18U  W=0.48U  
M13     u8_D    U22_in  VSS     VSS     N   L=0.18U  W=0.84U  
M14     u8_D    U22_in  VDD     VDD     P   L=0.18U  W=1.52U  
M15     U24_out u8_D    VSS     VSS     N   L=0.18U  W=0.72U  
M16     U24_out u8_D    VDD     VDD     P   L=0.185U  W=1.52U  
M17     u8_G    u8_GB   VSS     VSS     N   L=0.18U  W=0.47U  
M18     u8_G    u8_GB   VDD     VDD     P   L=0.186U  W=1.38U  
M19     u8_GB   CP      VSS     VSS     N   L=0.18U  W=0.69U  
M20     u8_GB   CP      VDD     VDD     P   L=0.18U  W=1.88U  
M21     U28_GB  U28_G   VSS     VSS     N   L=0.18U  W=0.62U  
M22     U28_GB  U28_G   VDD     VDD     P   L=0.185U  W=1.55U  
M23     U28_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M24     U28_D   D       VDD     VDD     P   L=0.185U  W=1.55U  
M25     U28_G   ENN     VSS     VSS     N   L=0.18U  W=0.62U  
M26     U28_G   ENN     VDD     VDD     P   L=0.185U  W=1.55U  
M27     u9_S    U23_in  VSS     VSS     N   L=0.18U  W=0.72U  
M28     u9_S    U23_in  VDD     VDD     P   L=0.186U  W=1.38U  
M29     Q       U23_in  VSS     VSS     N   L=0.182333U  W=2.91U  
M30     Q       U23_in  VDD     VDD     P   L=0.18U  W=8.2U  
M31     U27_D   u9_S    VSS     VSS     N   L=0.18U  W=0.62U  
M32     U27_D   u9_S    VDD     VDD     P   L=0.185U  W=1.52U  
M33     U23_in  u8_S    VSS     VSS     N   L=0.18U  W=0.92U  
M34     U23_in  u8_S    VDD     VDD     P   L=0.185U  W=1.66U  

.ENDS denrq4

.SUBCKT depfq4 Q  CPN D ENN SDN VDD VSS
M1      U32_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.83U  
M2      U32_out U32_in1 U32_u7_drain VSS     N   L=0.18U  W=0.83U  
M3      U32_out U32_in1 VDD     VDD     P   L=0.184U  W=1.58U  
M4      VDD     SDN     U32_out VDD     P   L=0.18U  W=1.25U  
M5      U35_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.75U  
M6      U35_out U35_in1 U35_u7_drain VSS     N   L=0.18U  W=0.75U  
M7      U35_out U35_in1 VDD     VDD     P   L=0.185U  W=1.59U  
M8      VDD     SDN     U35_out VDD     P   L=0.18U  W=1.59U  
M9      u8_S    u8_GB   U32_out VDD     P   L=0.187U  W=1.19U  
M10     u8_S    u8_G    U32_out VSS     N   L=0.18U  W=0.48U  
M11     U35_out u8_G    u8_S    VDD     P   L=0.187U  W=1.19U  
M12     U35_out u8_GB   u8_S    VSS     N   L=0.18U  W=0.48U  
M13     U24_out u8_GB   U32_in1 VDD     P   L=0.187U  W=1.11U  
M14     U24_out u8_G    U32_in1 VSS     N   L=0.18U  W=0.49U  
M15     U28_S   U30_out U28_D   VDD     P   L=0.185U  W=1.52U  
M16     U28_S   U30_in  U28_D   VSS     N   L=0.18U  W=0.62U  
M17     U32_in1 u8_G    U28_S   VDD     P   L=0.18U  W=1.11U  
M18     U32_in1 u8_GB   U28_S   VSS     N   L=0.18U  W=0.49U  
M19     U28_S   U30_in  U27_D   VDD     P   L=0.18U  W=1.45U  
M20     U28_S   U30_out U27_D   VSS     N   L=0.18U  W=0.62U  
M21     U24_out U32_out VSS     VSS     N   L=0.18U  W=0.65U  
M22     U24_out U32_out VDD     VDD     P   L=0.18U  W=1.3U  
M23     u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.48U  
M24     u8_GB   u8_G    VDD     VDD     P   L=0.18U  W=1.11U  
M25     u8_G    CPN     VSS     VSS     N   L=0.18U  W=0.69U  
M26     u8_G    CPN     VDD     VDD     P   L=0.184U  W=1.73U  
M27     U30_out U30_in  VSS     VSS     N   L=0.18U  W=0.62U  
M28     U30_out U30_in  VDD     VDD     P   L=0.18U  W=1.55U  
M29     U28_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M30     U28_D   D       VDD     VDD     P   L=0.18U  W=1.52U  
M31     U30_in  ENN     VSS     VSS     N   L=0.18U  W=0.62U  
M32     U30_in  ENN     VDD     VDD     P   L=0.185U  W=1.55U  
M33     Q       U35_in1 VSS     VSS     N   L=0.18U  W=2.91U  
M34     Q       U35_in1 VDD     VDD     P   L=0.182U  W=8.2U  
M35     U35_in1 u8_S    VSS     VSS     N   L=0.18U  W=0.69U  
M36     U35_in1 u8_S    VDD     VDD     P   L=0.185U  W=1.66U  
M37     U27_D   U35_out VSS     VSS     N   L=0.18U  W=0.62U  
M38     U27_D   U35_out VDD     VDD     P   L=0.186U  W=1.45U  

.ENDS depfq4

.SUBCKT deprq4 Q  CP D ENN SDN VDD VSS
M1      U32_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.83U  
M2      U32_out U32_in1 U32_u7_drain VSS     N   L=0.18U  W=0.83U  
M3      U32_out U32_in1 VDD     VDD     P   L=0.185U  W=1.56U  
M4      VDD     SDN     U32_out VDD     P   L=0.18U  W=1.14U  
M5      U35_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.83U  
M6      u9_S    U35_in1 U35_u7_drain VSS     N   L=0.18U  W=0.83U  
M7      u9_S    U35_in1 VDD     VDD     P   L=0.18U  W=1.63U  
M8      VDD     SDN     u9_S    VDD     P   L=0.185U  W=1.63U  
M9      u8_S    u8_GB   U32_out VDD     P   L=0.18U  W=1.11U  
M10     u8_S    u8_G    U32_out VSS     N   L=0.18U  W=0.48U  
M11     U24_out u8_GB   U32_in1 VDD     P   L=0.187U  W=1.11U  
M12     U24_out u8_G    U32_in1 VSS     N   L=0.18U  W=0.48U  
M13     u9_S    u8_G    u8_S    VDD     P   L=0.18U  W=1.11U  
M14     u9_S    u8_GB   u8_S    VSS     N   L=0.18U  W=0.48U  
M15     U28_S   U30_out U28_D   VDD     P   L=0.18U  W=1.52U  
M16     U28_S   U30_in  U28_D   VSS     N   L=0.18U  W=0.62U  
M17     U28_S   u8_G    U32_in1 VDD     P   L=0.18U  W=1.11U  
M18     U28_S   u8_GB   U32_in1 VSS     N   L=0.18U  W=0.48U  
M19     U28_S   U30_in  U27_D   VDD     P   L=0.185U  W=1.45U  
M20     U28_S   U30_out U27_D   VSS     N   L=0.18U  W=0.62U  
M21     U24_out U32_out VSS     VSS     N   L=0.18U  W=0.63U  
M22     U24_out U32_out VDD     VDD     P   L=0.18U  W=1.2U  
M23     u8_G    u8_GB   VSS     VSS     N   L=0.18U  W=0.48U  
M24     u8_G    u8_GB   VDD     VDD     P   L=0.187U  W=1.11U  
M25     u8_GB   CP      VSS     VSS     N   L=0.18U  W=0.69U  
M26     u8_GB   CP      VDD     VDD     P   L=0.184U  W=1.73U  
M27     U30_out U30_in  VSS     VSS     N   L=0.18U  W=0.62U  
M28     U30_out U30_in  VDD     VDD     P   L=0.18U  W=1.55U  
M29     U28_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M30     U28_D   D       VDD     VDD     P   L=0.185U  W=1.52U  
M31     U30_in  ENN     VSS     VSS     N   L=0.18U  W=0.62U  
M32     U30_in  ENN     VDD     VDD     P   L=0.185U  W=1.55U  
M33     Q       U35_in1 VSS     VSS     N   L=0.18U  W=2.77U  
M34     Q       U35_in1 VDD     VDD     P   L=0.183U  W=8.2U  
M35     U27_D   u9_S    VSS     VSS     N   L=0.18U  W=0.62U  
M36     U27_D   u9_S    VDD     VDD     P   L=0.18U  W=1.45U  
M37     U35_in1 u8_S    VSS     VSS     N   L=0.18U  W=0.69U  
M38     U35_in1 u8_S    VDD     VDD     P   L=0.185U  W=1.66U  

.ENDS deprq4

.SUBCKT dfbfb4 Q QN  CDN CPN D SDN VDD VSS
M1      u7_S    u7_GB   u7_D    VDD     P   L=0.187U   PD=.991U  W=1.25U
M2      u7_S    u7_G    u7_D    VSS     N   L=0.18U  PD=.850U  W=0.48U
M3      U19_out u7_G    u9_D    VDD     P   L=0.18U  PD=.914U  W=1.05U
M4      U19_out u7_GB   u9_D    VSS     N   L=0.18U    W=0.48U   
+  PD=1.370U
M5      U16_out u7_G    u7_D    VDD     P   L=0.18U    W=1.25U
M6      U16_out u7_GB   u7_D    VSS     N   L=0.18U    W=0.48U
M7      u14_in1 u7_GB   u9_D    VDD     P   L=0.18U   W=1.05U    
+  PD=1.086U
M8      u14_in1 u7_G    u9_D    VSS     N   L=0.18U   PD=.940U  W=0.48U
M9      U19_u7_drain SDN     VSS     VSS     N   L=0.18U    W=0.86U
+  PD=1.370U
M10     U19_out U19_in1 U19_u7_drain VSS     N   L=0.18U   W=0.86U
+  PS=1.370U PD=1.370U
M11     U19_out U19_in1 VDD     VDD     P   L=0.187U   W=1.25U
+  PD=.914U
M12     VDD     SDN     U19_out VDD     P   L=0.18U   PS=.914U  W=1.25U
M13     u14_u7_drain CDN     VSS     VSS     N   L=0.18U   W=0.87U
+  PD=.850U
M14     u7_S    u14_in1 u14_u7_drain VSS     N   L=0.18U   W=0.87U
+  PS=.850U PD=.850U
M15     u7_S    u14_in1 VDD     VDD     P   L=0.18U  PD=.991U  W=1.38U
M16     VDD     CDN     u7_S    VDD     P   L=0.186U  W=1.4U
+  PS=.991U
M17     u13_u7_drain SDN     VSS     VSS     N   L=0.18U   W=0.87U
+  PD=.940U
M18     u14_in1 u7_D    u13_u7_drain VSS     N   L=0.18U   W=0.87U
+  PS=.940U PD=.940U
M19     u14_in1 u7_D    VDD     VDD     P   L=0.189U    W=1.32U
+  PD=1.086U
M20     VDD     SDN     u14_in1 VDD     P   L=0.186U   W=1.32U
+  PS=1.086U
M21     u12_u7_drain CDN     VSS     VSS     N   L=0.18U     W=1U
+  PD=1.400U
M22     U19_in1 u9_D    u12_u7_drain VSS     N   L=0.18U    W=1U
+  PS=1.400U PD=1.400U
M23     U19_in1 u9_D    VDD     VDD     P   L=0.185U   W=1.52U
+  PD=1.305U
M24     VDD     CDN     U19_in1 VDD     P   L=0.187U   W=1.52U
+  PS=1.305U
M25     u7_G    CPN     VSS     VSS     N   L=0.18U    W=0.69U
M26     u7_G    CPN     VDD     VDD     P   L=0.18U   W=1.73U
M27     u7_GB   u7_G    VSS     VSS     N   L=0.18U   W=0.55U
M28     u7_GB   u7_G    VDD     VDD     P   L=0.187U   W=1.52U
M29     U16_out D       VSS     VSS     N   L=0.18U   W=0.62U
M30     U16_out D       VDD     VDD     P   L=0.186U     W=1.45U
M31     Q       U19_in1 VSS     VSS     N   L=0.18U    W=2.95U
M32     Q       U19_in1 VDD     VDD     P   L=0.182U    W=8.2U
M33     QN      u9_D    VSS     VSS     N   L=0.18U   W=2.82U
M34     QN      u9_D    VDD     VDD     P   L=0.182U   W=8.34U

.ENDS dfbfb4

.SUBCKT dfbrb4 Q QN  CDN CP D SDN VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.18U  W=1.11U   
+  PS=1.053U
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U  W=0.48U   PS=.900U
M3      U15_S   u8_G    U15_D   VDD     P   L=0.18U  W=1.25U  
M4      U15_S   u8_GB   U15_D   VSS     N   L=0.18U  W=0.48U  
M5      u7_S    u8_GB   U15_S   VDD     P   L=0.18U  W=1.11U   PD=.940U
M6      u7_S    u8_G    U15_S   VSS     N   L=0.18U  W=0.48U   PD=.855U
M7      U24_out u8_G    u8_S    VDD     P   L=0.18U  W=1.11U   
+  PD=1.155U
M8      U24_out u8_GB   u8_S    VSS     N   L=0.18U  W=0.48U   PD=.755U
M9      u8_G    u8_GB   VSS     VSS     N   L=0.18U  W=0.55U  
M10     u8_G    u8_GB   VDD     VDD     P   L=0.18U  W=1.52U  
M11     u8_GB   CP      VSS     VSS     N   L=0.18U  W=0.69U  
M12     u8_GB   CP      VDD     VDD     P   L=0.184U  W=1.73U  
M13     U15_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M14     U15_D   D       VDD     VDD     P   L=0.186U  W=1.45U  
M15     Q       U24_in1 VSS     VSS     N   L=0.18U  W=2.89U  
M16     Q       U24_in1 VDD     VDD     P   L=0.18225U  W=8.2U  
M17     QN      u8_S    VSS     VSS     N   L=0.18U  W=2.89U  
M18     QN      u8_S    VDD     VDD     P   L=0.182U  W=8.2U  
M19     U21_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.87U   
+  PD=.900U
M20     u8_D    U15_S   U21_u7_drain VSS     N   L=0.18U  W=0.87U   
+  PS=.900U PD=.900U
M21     u8_D    U15_S   VDD     VDD     P   L=0.186U  W=1.32U   
+  PD=1.053U
M22     VDD     SDN     u8_D    VDD     P   L=0.186U  W=1.32U   
+  PS=1.053U
M23     U22_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.87U   
+  PD=.855U
M24     u7_S    u8_D    U22_u7_drain VSS     N   L=0.18U  W=0.94U   
+  PS=.855U PD=.855U
M25     u7_S    u8_D    VDD     VDD     P   L=0.186U  W=1.38U   PD=.940U
M26     VDD     CDN     u7_S    VDD     P   L=0.186U  W=1.38U   
+  PS=.940U
M27     U24_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.91U   
+  PD=.755U
M28     U24_out U24_in1 U24_u7_drain VSS     N   L=0.18U  W=0.91U   
+  PS=.755U PD=.755U
M29     U24_out U24_in1 VDD     VDD     P   L=0.187U  W=1.25U   
+  PD=1.155U
M30     VDD     SDN     U24_out VDD     P   L=0.187U  W=1.25U   
+  PS=1.155U
M31     U23_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.96U   
+  PD=1.027U
M32     U24_in1 u8_S    U23_u7_drain VSS     N   L=0.18U  W=0.96U   
+  PS=1.027U PD=1.065U
M33     U24_in1 u8_S    VDD     VDD     P   L=0.18U  W=1.52U   
+  PD=1.437U
M34     VDD     CDN     U24_in1 VDD     P   L=0.185U  W=1.52U   
+  PS=1.437U

.ENDS dfbrb4

.SUBCKT dfcfb4 Q QN  CDN CPN D VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.18U  W=1.14U  
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U  W=0.66U  
M3      u7_S    u8_GB   u7_D    VDD     P   L=0.189U  W=1.25U   PD=.921U
M4      u7_S    u8_G    u7_D    VSS     N   L=0.18U  W=0.48U   PD=.750U
M5      u7_D    u8_G    U15_D   VDD     P   L=0.186U  W=1.25U  
M6      u7_D    u8_GB   U15_D   VSS     N   L=0.18U  W=0.48U  
M7      U23_out u8_G    u8_S    VDD     P   L=0.187U  W=1.14U  
M8      U23_out u8_GB   u8_S    VSS     N   L=0.18U  W=0.55U  
M9      u8_G    CPN     VSS     VSS     N   L=0.18U  W=0.69U  
M10     u8_G    CPN     VDD     VDD     P   L=0.185U  W=1.73U  
M11     u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.55U  
M12     u8_GB   u8_G    VDD     VDD     P   L=0.18U  W=1.52U  
M13     U15_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M14     U15_D   D       VDD     VDD     P   L=0.18U  W=1.45U  
M15     u8_D    u7_D    VSS     VSS     N   L=0.18U  W=0.64U  
M16     u8_D    u7_D    VDD     VDD     P   L=0.185U  W=1.43U  
M17     U23_out U24_out VSS     VSS     N   L=0.18U  W=0.47U  
M18     U23_out U24_out VDD     VDD     P   L=0.18U  W=1.02U  
M19     Q       U24_out VSS     VSS     N   L=0.18U  W=2.88U  
M20     Q       U24_out VDD     VDD     P   L=0.1836U  W=8.2U  
M21     QN      u8_S    VSS     VSS     N   L=0.18U  W=2.88U  
M22     QN      u8_S    VDD     VDD     P   L=0.1832U  W=8.2U  
M23     U25_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.87U   
+  PD=.750U
M24     u7_S    u8_D    U25_u7_drain VSS     N   L=0.18U  W=0.87U   
+  PS=.750U PD=.750U
M25     u7_S    u8_D    VDD     VDD     P   L=0.185U  W=1.52U   
+  PD=.921U
M26     VDD     CDN     u7_S    VDD     P   L=0.185U  W=1.52U   PS=.921U
M27     U24_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.86U   
+  PD=1.045U
M28     U24_out u8_S    U24_u7_drain VSS     N   L=0.18U  W=0.86U   
+  PS=1.045U PD=1.045U
M29     U24_out u8_S    VDD     VDD     P   L=0.18U  W=1.63U   
+  PD=1.094U
M30     VDD     CDN     U24_out VDD     P   L=0.184U  W=1.63U   
+  PS=1.094U

.ENDS dfcfb4

.SUBCKT dfcfq4 Q  CDN CPN D VDD VSS
M1      U25_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.87U   
+  PD=.750U
M2      U25_out U25_in1 U25_u7_drain VSS     N   L=0.18U  W=0.87U   
+  PS=.750U PD=.750U
M3      U25_out U25_in1 VDD     VDD     P   L=0.185U  W=1.52U   PD=.939U
M4      VDD     CDN     U25_out VDD     P   L=0.18U  W=1.52U   
+  PS=.939U
M5      U24_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.86U   
+  PD=1.575U
M6      U24_out U24_in1 U24_u7_drain VSS     N   L=0.18U  W=0.86U   
+  PS=1.575U PD=1.575U
M7      U24_out U24_in1 VDD     VDD     P   L=0.185U  W=1.63U   
+  PD=1.175U
M8      VDD     CDN     U24_out VDD     P   L=0.18U  W=1.63U   
+  PS=1.175U
M9      U25_in1 U22_in  VSS     VSS     N   L=0.18U  W=0.64U  
M10     U25_in1 U22_in  VDD     VDD     P   L=0.18U  W=1.43U  
M11     u10_out CPN     VSS     VSS     N   L=0.18U  W=0.69U  
M12     u10_out CPN     VDD     VDD     P   L=0.184U  W=1.73U  
M13     u11_out u10_out VSS     VSS     N   L=0.18U  W=0.55U  
M14     u11_out u10_out VDD     VDD     P   L=0.18U  W=1.52U  
M15     U15_S   D       VSS     VSS     N   L=0.18U  W=0.62U  
M16     U15_S   D       VDD     VDD     P   L=0.18U  W=1.45U  
M17     U23_out U24_out VSS     VSS     N   L=0.18U  W=0.47U  
M18     U23_out U24_out VDD     VDD     P   L=0.18U  W=1.02U  
M19     Q       U24_out VSS     VSS     N   L=0.1825U  W=2.85U  
M20     Q       U24_out VDD     VDD     P   L=0.182U  W=8.32U  
M21     U15_S   u10_out U22_in  VDD     P   L=0.186U  W=1.25U  
M22     U15_S   u11_out U22_in  VSS     N   L=0.18U  W=0.48U  
M23     U22_in  u11_out U25_out VDD     P   L=0.18U  W=1.25U   PS=.939U
M24     U22_in  u10_out U25_out VSS     N   L=0.18U  W=0.48U   PS=.750U
M25     U24_in1 u10_out U23_out VDD     P   L=0.187U  W=1.14U  
M26     U24_in1 u11_out U23_out VSS     N   L=0.18U  W=0.55U  
M27     U25_in1 u11_out U24_in1 VDD     P   L=0.187U  W=1.14U  
M28     U25_in1 u10_out U24_in1 VSS     N   L=0.18U  W=0.66U  

.ENDS dfcfq4

.SUBCKT dfcrb4 Q QN  CDN CP D VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.18U  W=1.14U  
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U  W=0.66U  
M3      u7_S    u8_GB   u7_D    VDD     P   L=0.18U  W=1.25U   
+  PD=1.078U
M4      u7_S    u8_G    u7_D    VSS     N   L=0.18U  W=0.48U   PD=.750U
M5      u7_D    u8_G    U15_D   VDD     P   L=0.187U  W=1.25U  
M6      u7_D    u8_GB   U15_D   VSS     N   L=0.18U  W=0.48U  
M7      U23_out u8_G    u8_S    VDD     P   L=0.187U  W=1.14U  
M8      U23_out u8_GB   u8_S    VSS     N   L=0.18U  W=0.55U  
M9      u8_G    u8_GB   VSS     VSS     N   L=0.18U  W=0.55U  
M10     u8_G    u8_GB   VDD     VDD     P   L=0.18U  W=1.52U  
M11     u8_GB   CP      VSS     VSS     N   L=0.18U  W=0.69U  
M12     u8_GB   CP      VDD     VDD     P   L=0.185U  W=1.73U  
M13     u8_D    u7_D    VSS     VSS     N   L=0.18U  W=0.64U  
M14     u8_D    u7_D    VDD     VDD     P   L=0.186U  W=1.43U  
M15     U15_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M16     U15_D   D       VDD     VDD     P   L=0.18U  W=1.45U  
M17     U23_out U24_out VSS     VSS     N   L=0.18U  W=0.47U  
M18     U23_out U24_out VDD     VDD     P   L=0.18U  W=1.02U  
M19     QN      u8_S    VSS     VSS     N   L=0.18U  W=2.91U  
M20     QN      u8_S    VDD     VDD     P   L=0.182U  W=8.2U  
M21     Q       U24_out VSS     VSS     N   L=0.18U  W=2.91U  
M22     Q       U24_out VDD     VDD     P   L=0.182U  W=8.2U  
M23     U25_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.87U   
+  PD=.750U
M24     u7_S    u8_D    U25_u7_drain VSS     N   L=0.18U  W=0.87U   
+  PS=.750U PD=.750U
M25     u7_S    u8_D    VDD     VDD     P   L=0.185U  W=1.52U   
+  PD=1.078U
M26     VDD     CDN     u7_S    VDD     P   L=0.185U  W=1.52U   
+  PS=1.078U
M27     U24_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.86U   
+  PD=1.045U
M28     U24_out u8_S    U24_u7_drain VSS     N   L=0.18U  W=0.86U   
+  PS=1.045U PD=1.045U
M29     U24_out u8_S    VDD     VDD     P   L=0.18U  W=1.63U   
+  PD=1.079U
M30     VDD     CDN     U24_out VDD     P   L=0.185U  W=1.63U   
+  PS=1.079U

.ENDS dfcrb4

.SUBCKT dfcrn4 QN  CDN CP D VDD VSS
M1      U25_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.87U   
+  PD=.785U
M2      U25_out U25_in1 U25_u7_drain VSS     N   L=0.18U  W=0.87U   
+  PS=.785U PD=.785U
M3      U25_out U25_in1 VDD     VDD     P   L=0.185U  W=1.52U   
+  PD=1.130U
M4      VDD     CDN     U25_out VDD     P   L=0.18U  W=1.52U   
+  PS=1.130U
M5      U24_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.86U   
+  PD=.750U
M6      U24_out u9_D    U24_u7_drain VSS     N   L=0.18U  W=0.86U   
+  PS=.750U PD=.750U
M7      U24_out u9_D    VDD     VDD     P   L=0.18U  W=1.63U   PD=.790U
M8      VDD     CDN     U24_out VDD     P   L=0.185U  W=1.63U   PS=.790U
M9      U25_in1 U22_in  VSS     VSS     N   L=0.18U  W=0.64U  
M10     U25_in1 U22_in  VDD     VDD     P   L=0.18U  W=1.43U  
M11     u10_out CP      VSS     VSS     N   L=0.18U  W=0.69U  
M12     u10_out CP      VDD     VDD     P   L=0.184U  W=1.73U  
M13     u11_out u10_out VSS     VSS     N   L=0.18U  W=0.55U  
M14     u11_out u10_out VDD     VDD     P   L=0.18U  W=1.52U  
M15     U15_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M16     U15_D   D       VDD     VDD     P   L=0.18U  W=1.45U  
M17     QN      u9_D    VSS     VSS     N   L=0.18U  W=2.89U  
M18     QN      u9_D    VDD     VDD     P   L=0.1825U  W=8.2U  
M19     u9_S    U24_out VSS     VSS     N   L=0.18U  W=0.47U  
M20     u9_S    U24_out VDD     VDD     P   L=0.18U  W=1.02U  
M21     U25_out u10_out U22_in  VDD     P   L=0.18U  W=1.25U   
+  PD=1.130U
M22     U25_out u11_out U22_in  VSS     N   L=0.18U  W=0.48U   PD=.785U
M23     U22_in  u11_out U15_D   VDD     P   L=0.187U  W=1.25U  
M24     U22_in  u10_out U15_D   VSS     N   L=0.18U  W=0.48U  
M25     u9_S    u11_out u9_D    VDD     P   L=0.18U  W=1.14U  
M26     u9_S    u10_out u9_D    VSS     N   L=0.18U  W=0.55U  
M27     U25_in1 u10_out u9_D    VDD     P   L=0.187U  W=1.14U  
M28     U25_in1 u11_out u9_D    VSS     N   L=0.18U  W=0.66U  

.ENDS dfcrn4

.SUBCKT dfcrq4 CP CDN D Q VDD VSS 
M1      u8_S    u8_GB   u8_D    VDD     P   L=.1800U  W=1.1400U  
M2      u8_S    u8_G    u8_D    VSS     N   L=.1800U  W=.6600U  
M3      u7_S    u8_GB   U22_in  VDD     P   L=.1850U  W=1.2500U  
M4      u7_S    u8_G    U22_in  VSS     N   L=.1800U  W=.4800U  
M5      U15_S   u8_G    U22_in  VDD     P   L=.1850U  W=1.2500U  
M6      U15_S   u8_GB   U22_in  VSS     N   L=.1800U  W=.4800U  
M7      U23_out u8_G    u8_S    VDD     P   L=.1860U  W=1.1400U  
M8      U23_out u8_GB   u8_S    VSS     N   L=.1800U  W=.5500U  
M9      u8_D    U22_in  VSS     VSS     N   L=.1800U  W=.6400U  
M10     u8_D    U22_in  VDD     VDD     P   L=.1850U  W=1.4200U  
M11     u8_GB   CP      VSS     VSS     N   L=.1800U  W=.6900U  
M12     u8_GB   CP      VDD     VDD     P   L=.1840U  W=1.7300U  
M13     u8_G    u8_GB   VSS     VSS     N   L=.1800U  W=.5500U  
M14     u8_G    u8_GB   VDD     VDD     P   L=.1800U  W=1.5200U  
M15     U15_S   D       VSS     VSS     N   L=.1800U  W=.6200U  
M16     U15_S   D       VDD     VDD     P   L=.1850U  W=1.4500U  
M17     U23_out U24_out VSS     VSS     N   L=.1800U  W=.4700U  
M18     U23_out U24_out VDD     VDD     P   L=.1870U  W=1.0200U  
M19     Q       U24_out VSS     VSS     N   L=.1800U  W=2.8900U  
M20     Q       U24_out VDD     VDD     P   L=.1840U  W=8.4000U  
M21     U25_u7_drain CDN     VSS     VSS     N   L=.1800U  W=.8700U  
M22     u7_S    u8_D    U25_u7_drain VSS     N   L=.1800U  W=.8700U  
M23     u7_S    u8_D    VDD     VDD     P   L=.1800U  W=1.5200U  
M24     VDD     CDN     u7_S    VDD     P   L=.1840U  W=1.5200U  
M25     U24_u7_drain CDN     VSS     VSS     N   L=.1800U  W=.8600U  
M26     U24_out u8_S    U24_u7_drain VSS     N   L=.1800U  W=.8600U  
M27     U24_out u8_S    VDD     VDD     P   L=.1840U  W=1.6300U  
M28     VDD     CDN     U24_out VDD     P   L=.1800U  W=1.6300U  

.ENDS dfcrq4

.SUBCKT dfnfb4 Q QN  CPN D VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.18U  W=1.14U  
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U  W=0.64U  
M3      U24_out u8_GB   u7_D    VDD     P   L=0.189U  W=1.25U  
M4      U24_out u8_G    u7_D    VSS     N   L=0.18U  W=0.48U  
M5      u7_D    u8_G    U15_D   VDD     P   L=0.18U  W=1.25U  
M6      u7_D    u8_GB   U15_D   VSS     N   L=0.18U  W=0.48U  
M7      u9_S    u8_G    u8_S    VDD     P   L=0.18U  W=1.14U  
M8      u9_S    u8_GB   u8_S    VSS     N   L=0.18U  W=0.55U  
M9      U24_out u8_D    VSS     VSS     N   L=0.18U  W=0.86U  
M10     U24_out u8_D    VDD     VDD     P   L=0.18U  W=1.74U  
M11     u8_G    CPN     VSS     VSS     N   L=0.18U  W=0.69U  
M12     u8_G    CPN     VDD     VDD     P   L=0.184U  W=1.73U  
M13     u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.55U  
M14     u8_GB   u8_G    VDD     VDD     P   L=0.18U  W=1.52U  
M15     u8_D    u7_D    VSS     VSS     N   L=0.18U  W=0.72U  
M16     u8_D    u7_D    VDD     VDD     P   L=0.185U  W=1.74U  
M17     U15_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M18     U15_D   D       VDD     VDD     P   L=0.185U  W=1.45U  
M19     u9_S    U23_in  VSS     VSS     N   L=0.18U  W=0.72U  
M20     u9_S    U23_in  VDD     VDD     P   L=0.184U  W=1.88U  
M21     QN      u8_S    VSS     VSS     N   L=0.18U  W=2.89U  
M22     QN      u8_S    VDD     VDD     P   L=0.18U  W=8.25U  
M23     Q       U23_in  VSS     VSS     N   L=0.182U  W=2.89U  
M24     Q       U23_in  VDD     VDD     P   L=0.184U  W=8.21U  
M25     U23_in  u8_S    VSS     VSS     N   L=0.18U  W=.83U  
M26     U23_in  u8_S    VDD     VDD     P   L=0.184U  W=1.88U  

.ENDS dfnfb4

.SUBCKT dfnrb4 Q QN  CP D VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.187U  W=1.14U  
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U   W=0.64U  
M3      u7_S    u8_GB   u7_D    VDD     P   L=0.18U   W=1.25U  
M4      u7_S    u8_G    u7_D    VSS     N   L=0.18U   W=0.48U  
M5      u7_D    u8_G    U15_D   VDD     P   L=0.187U  W=1.25U  
M6      u7_D    u8_GB   U15_D   VSS     N   L=0.18U   W=0.48U  
M7      U23_out u8_G    u8_S    VDD     P   L=0.18U   W=1.14U  
M8      U23_out u8_GB   u8_S    VSS     N   L=0.18U   W=0.55U  
M9      u8_GB   CP      VSS     VSS     N   L=0.18U   W=0.69U  
M10     u8_GB   CP      VDD     VDD     P   L=0.184U   W=1.73U  
M11     u8_G    u8_GB   VSS     VSS     N   L=0.18U   W=0.55U  
M12     u8_G    u8_GB   VDD     VDD     P   L=0.18U   W=1.52U  
M13     U15_D   D       VSS     VSS     N   L=0.18U   W=0.62U  
M14     U15_D   D       VDD     VDD     P   L=0.18U   W=1.45U  
M15     u8_D    u7_D    VSS     VSS     N   L=0.18U   W=0.72U  
M16     u8_D    u7_D    VDD     VDD     P   L=0.18U   W=1.74U  
M17     u7_S    u8_D    VSS     VSS     N   L=0.18U   W=0.86U  
M18     u7_S    u8_D    VDD     VDD     P   L=0.185U  W=1.74U  
M19     U23_out U23_in  VSS     VSS     N   L=0.18U   W=0.72U  
M20     U23_out U23_in  VDD     VDD     P   L=0.184U  W=1.88U  
M21     U23_in  u8_S    VSS     VSS     N   L=0.18U   W=0.83U
M22     U23_in  u8_S    VDD     VDD     P   L=0.18U   W=1.88U  
M23     Q       U23_in  VSS     VSS     N   L=0.18U   W=2.89U  
M24     Q       U23_in  VDD     VDD     P   L=0.182U  W=8.2U  
M25     QN      u8_S    VSS     VSS     N   L=0.18U   W=2.89U  
M26     QN      u8_S    VDD     VDD     P   L=0.182U  W=8.2U  

.ENDS dfnrb4

.SUBCKT dfnrn4 QN  CP D VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.187U  W=1.14U  
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U  W=0.64U  
M3      U15_S   u8_G    U15_D   VDD     P   L=0.18U  W=1.25U  
M4      U15_S   u8_GB   U15_D   VSS     N   L=0.18U  W=0.48U  
M5      u7_S    u8_GB   U15_S   VDD     P   L=0.187U  W=1.25U  
M6      u7_S    u8_G    U15_S   VSS     N   L=0.18U  W=0.48U  
M7      U23_out u8_G    u8_S    VDD     P   L=0.18U  W=1.14U  
M8      U23_out u8_GB   u8_S    VSS     N   L=0.18U  W=0.55U  
M9      u8_GB   CP      VSS     VSS     N   L=0.18U  W=0.69U  
M10     u8_GB   CP      VDD     VDD     P   L=0.184U  W=1.73U  
M11     u8_G    u8_GB   VSS     VSS     N   L=0.18U  W=0.55U  
M12     u8_G    u8_GB   VDD     VDD     P   L=0.185U  W=1.52U  
M13     u8_D    U15_S   VSS     VSS     N   L=0.18U  W=0.72U  
M14     u8_D    U15_S   VDD     VDD     P   L=0.184U  W=1.74U  
M15     U15_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M16     U15_D   D       VDD     VDD     P   L=0.186U  W=1.45U  
M17     u7_S    u8_D    VSS     VSS     N   L=0.18U  W=0.86U  
M18     u7_S    u8_D    VDD     VDD     P   L=0.185U  W=1.74U  
M19     U25_out u8_S    VSS     VSS     N   L=0.18U  W=0.83U  
M20     U25_out u8_S    VDD     VDD     P   L=0.184U  W=1.87U  
M21     U23_out U25_out VSS     VSS     N   L=0.18U  W=0.72U  
M22     U23_out U25_out VDD     VDD     P   L=0.184U  W=1.87U  
M23     QN      u8_S    VSS     VSS     N   L=0.18U  W=2.89U  
M24     QN      u8_S    VDD     VDD     P   L=0.184U  W=8.4U  

.ENDS dfnrn4

.SUBCKT dfnrq4 Q  CP D VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.18U  W=1.14U  
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U  W=0.64U  
M3      U22_in  u8_G    U15_D   VDD     P   L=0.18U  W=1.25U  
M4      U22_in  u8_GB   U15_D   VSS     N   L=0.18U  W=0.48U  
M5      U24_out u8_GB   U22_in  VDD     P   L=0.186U  W=1.25U  
M6      U24_out u8_G    U22_in  VSS     N   L=0.18U  W=0.48U  
M7      u9_S    u8_G    u8_S    VDD     P   L=0.187U  W=1.14U  
M8      u9_S    u8_GB   u8_S    VSS     N   L=0.18U  W=0.55U  
M9      u8_D    U22_in  VSS     VSS     N   L=0.18U  W=0.72U  
M10     u8_D    U22_in  VDD     VDD     P   L=0.18U  W=1.74U  
M11     U24_out u8_D    VSS     VSS     N   L=0.18U  W=0.86U  
M12     U24_out u8_D    VDD     VDD     P   L=0.185U  W=1.74U  
M13     u8_GB   CP      VSS     VSS     N   L=0.18U  W=0.69U  
M14     u8_GB   CP      VDD     VDD     P   L=0.185U  W=1.73U  
M15     u8_G    u8_GB   VSS     VSS     N   L=0.18U  W=0.55U  
M16     u8_G    u8_GB   VDD     VDD     P   L=0.18U  W=1.52U  
M17     U15_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M18     U15_D   D       VDD     VDD     P   L=0.186U  W=1.45U  
M19     Q       u3_in   VSS     VSS     N   L=0.18U  W=2.89U  
M20     Q       u3_in   VDD     VDD     P   L=0.183U  W=8.4U  
M21     u3_in   u8_S    VSS     VSS     N   L=0.18U  W=0.83U  
M22     u3_in   u8_S    VDD     VDD     P   L=0.18U  W=1.87U  
M23     u9_S    u3_in   VSS     VSS     N   L=0.18U  W=0.72U  
M24     u9_S    u3_in   VDD     VDD     P   L=0.184U  W=1.87U  

.ENDS dfnrq4

.SUBCKT dfpfb4 Q QN  CPN D SDN VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.18U  W=1.05U   
+  PS=1.036U
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U  W=0.48U   PS=.990U
M3      u7_S    u8_GB   u7_D    VDD     P   L=0.18U  W=1.25U  
M4      u7_S    u8_G    u7_D    VSS     N   L=0.18U  W=0.48U  
M5      u7_D    u8_G    U15_D   VDD     P   L=0.186U  W=1.25U  
M6      u7_D    u8_GB   U15_D   VSS     N   L=0.18U  W=0.48U  
M7      U24_out u8_G    u8_S    VDD     P   L=0.18U  W=1.05U   
+  PD=1.102U
M8      U24_out u8_GB   u8_S    VSS     N   L=0.18U  W=0.48U   PD=.705U
M9      u8_G    CPN     VSS     VSS     N   L=0.18U  W=0.69U  
M10     u8_G    CPN     VDD     VDD     P   L=0.185U  W=1.73U  
M11     u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.55U  
M12     u8_GB   u8_G    VDD     VDD     P   L=0.18U  W=1.52U  
M13     U15_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M14     U15_D   D       VDD     VDD     P   L=0.18U  W=1.45U  
M15     u7_S    u8_D    VSS     VSS     N   L=0.18U  W=0.87U  
M16     u7_S    u8_D    VDD     VDD     P   L=0.186U  W=1.45U  
M17     U24_in1 u8_S    VSS     VSS     N   L=0.18U  W=0.86U  
M18     U24_in1 u8_S    VDD     VDD     P   L=0.18U  W=1.87U  
M19     Q       U24_in1 VSS     VSS     N   L=0.18U  W=2.92U  
M20     Q       U24_in1 VDD     VDD     P   L=0.182U  W=8.2U  
M21     QN      u8_S    VSS     VSS     N   L=0.18U  W=2.92U  
M22     QN      u8_S    VDD     VDD     P   L=0.182U  W=8.2U  
M23     U25_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.87U   
+  PD=.990U
M24     u8_D    u7_D    U25_u7_drain VSS     N   L=0.18U  W=0.87U   
+  PS=.990U PD=.990U
M25     u8_D    u7_D    VDD     VDD     P   L=0.186U  W=1.32U   
+  PD=1.036U
M26     VDD     SDN     u8_D    VDD     P   L=0.186U  W=1.32U   
+  PS=1.036U
M27     U24_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.86U   
+  PD=.705U
M28     U24_out U24_in1 U24_u7_drain VSS     N   L=0.18U  W=0.86U   
+  PS=.705U PD=.705U
M29     U24_out U24_in1 VDD     VDD     P   L=0.186U  W=1.23U   
+  PD=1.102U
M30     VDD     SDN     U24_out VDD     P   L=0.18U  W=1.23U   
+  PS=1.102U

.ENDS dfpfb4

.SUBCKT dfprb4 Q QN  CP D SDN VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.186U  W=1.05U   
+  PS=1.173U
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U  W=0.48U   PS=.990U
M3      U15_S   u8_G    U15_D   VDD     P   L=0.187U  W=1.25U  
M4      U15_S   u8_GB   U15_D   VSS     N   L=0.18U  W=0.48U  
M5      u7_S    u8_GB   U15_S   VDD     P   L=0.18U  W=1.25U  
M6      u7_S    u8_G    U15_S   VSS     N   L=0.18U  W=0.48U  
M7      U24_out u8_G    u8_S    VDD     P   L=0.18U  W=1.05U   
+  PD=1.140U
M8      U24_out u8_GB   u8_S    VSS     N   L=0.18U  W=0.48U   PD=.770U
M9      u8_GB   CP      VSS     VSS     N   L=0.18U  W=0.69U  
M10     u8_GB   CP      VDD     VDD     P   L=0.184U  W=1.73U  
M11     u8_G    u8_GB   VSS     VSS     N   L=0.18U  W=0.55U  
M12     u8_G    u8_GB   VDD     VDD     P   L=0.18U  W=1.52U  
M13     U15_D   D       VSS     VSS     N   L=0.18U  W=0.62U  
M14     U15_D   D       VDD     VDD     P   L=0.18U  W=1.45U  
M15     u7_S    u8_D    VSS     VSS     N   L=0.18U  W=0.87U  
M16     u7_S    u8_D    VDD     VDD     P   L=0.186U  W=1.45U  
M17     U24_in1 u8_S    VSS     VSS     N   L=0.18U  W=0.86U  
M18     U24_in1 u8_S    VDD     VDD     P   L=0.18U  W=1.87U  
M19     Q       U24_in1 VSS     VSS     N   L=0.18U  W=2.92U  
M20     Q       U24_in1 VDD     VDD     P   L=0.18225U  W=8.2U  
M21     QN      u8_S    VSS     VSS     N   L=0.18U  W=2.92U  
M22     QN      u8_S    VDD     VDD     P   L=0.18U  W=8.2U  
M23     U25_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.87U   
+  PD=.990U
M24     u8_D    U15_S   U25_u7_drain VSS     N   L=0.18U  W=0.87U   
+  PS=.990U PD=.990U
M25     u8_D    U15_S   VDD     VDD     P   L=0.18U  W=1.32U   
+  PD=1.173U
M26     VDD     SDN     u8_D    VDD     P   L=0.186U  W=1.32U   
+  PS=1.173U
M27     U24_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.86U   
+  PD=.770U
M28     U24_out U24_in1 U24_u7_drain VSS     N   L=0.18U  W=0.86U   
+  PS=.770U PD=.770U
M29     U24_out U24_in1 VDD     VDD     P   L=0.186U  W=1.23U   
+  PD=1.140U
M30     VDD     SDN     U24_out VDD     P   L=0.18U  W=1.23U   
+  PS=1.140U

.ENDS dfprb4

.SUBCKT dl01d2 Z  I VDD VSS
M1      U65_drain U65_gate VDD     VDD     P   L=0.33U  W=0.44U
M2      U65_gate U79_gate VDD     VDD     P   L=0.3U  W=0.33U
M3      U79_gate I       VDD     VDD     P   L=0.184U  W=1.84U
M4      Z       U65_drain VDD     VDD     P   L=0.182U  W=4.1U
M5      U65_gate U79_gate VSS     VSS     N   L=0.18U  W=0.24U
M6      U65_drain U65_gate VSS     VSS     N   L=0.44U  W=0.25U
M7      U79_gate I       VSS     VSS     N   L=0.18U  W=0.42U
M8      Z       U65_drain VSS     VSS     N   L=0.18U  W=1.38U

.ENDS dl01d2

.SUBCKT dl01d4 Z  I VDD VSS
M1      U65_drain U65_gate VDD     VDD     P   L=0.21U  W=0.48U  
M2      U65_gate U79_gate VDD     VDD     P   L=0.19U  W=0.36U  
M3      U79_gate I       VDD     VDD     P   L=0.184U  W=1.92U  
M4      Z       U65_drain VDD     VDD     P   L=0.183U  W=8.2U  
M5      U65_gate U79_gate VSS     VSS     N   L=0.19U  W=0.24U  
M6      U65_drain U65_gate VSS     VSS     N   L=0.42U  W=0.36U  
M7      U79_gate I       VSS     VSS     N   L=0.18U  W=0.5U  
M8      Z       U65_drain VSS     VSS     N   L=0.185U  W=2.95U  

.ENDS dl01d4

.SUBCKT dl02d2 Z  I VDD VSS
M1      U65_drain U65_gate VDD     VDD     P   L=0.48U    W=0.34U
M2      U65_gate U79_gate VDD     VDD     P   L=0.9U    W=0.33U
M3      U79_gate I       VDD     VDD     P   L=0.184U     W=1.84U
M4      Z       U65_drain VDD     VDD     P   L=0.184U    W=4.10U
M5      U65_gate U79_gate VSS     VSS     N   L=0.83U     W=0.24U
M6      U65_drain U65_gate VSS     VSS     N   L=0.45U     W=0.24U
M7      U79_gate I       VSS     VSS     N   L=0.180U     W=0.42U
M8      Z       U65_drain VSS     VSS     N   L=0.180U     W=1.39U

.ENDS dl02d2

.SUBCKT dl02d4 Z  I VDD VSS
M1      U65_drain U65_gate VDD     VDD     P   L=0.34U    W=0.34U
M2      U65_gate U79_gate VDD     VDD     P   L=0.7U       W=0.33U
M3      U79_gate I       VDD     VDD     P   L=0.184U       W=1.84U
M4      Z       U65_drain VDD     VDD     P   L=0.183U      W=8.2U
M5      U65_gate U79_gate VSS     VSS     N   L=0.47U      W=0.24U
M6      U65_drain U65_gate VSS     VSS     N   L=0.5U    W=0.24U
M7      U79_gate I       VSS     VSS     N   L=0.18U       W=0.42U
M8      Z       U65_drain VSS     VSS     N   L=0.18U      W=2.77U

.ENDS dl02d4

.SUBCKT dl03d2 Z  I VDD VSS
M1      U8_drain U8_gate VDD     VDD     P   L=0.47U  W=0.42U
M2      U8_gate U6_gate VDD     VDD     P   L=1.66U  W=0.42U
M3      U1_drain I       VDD     VDD     P   L=0.184U  W=1.94U
M4      U6_gate U1_drain VDD     VDD     P   L=1.0U  W=0.42U
M5      Z       U9_drain VDD     VDD     P   L=0.184U  W=4.1U
M6      U9_drain U8_drain VDD     VDD     P   L=0.18U  W=0.42U
M7      U8_drain U8_gate VSS     VSS     N   L=0.75U  W=0.24U
M8      U8_gate U6_gate VSS     VSS     N   L=1.3U  W=0.24U
M9      U1_drain I       VSS     VSS     N   L=0.18U  W=0.42U
M10     U6_gate U1_drain VSS     VSS     N   L=0.95U  W=0.24U
M11     U9_drain U8_drain VSS     VSS     N   L=0.18U  W=0.44U
M12     Z       U9_drain VSS     VSS     N   L=0.189U  W=1.65U

.ENDS dl03d2

.SUBCKT dl03d4 Z  I VDD VSS
M1      U8_drain U8_gate VDD     VDD     P   L=0.42U  W=0.42U
M2      U8_gate U6_gate VDD     VDD     P   L=1.52U  W=0.42U
M3      U1_drain I       VDD     VDD     P   L=0.184U  W=1.94U
M4      U6_gate U1_drain VDD     VDD     P   L=0.97U  W=0.42U
M5      Z       U9_drain VDD     VDD     P   L=0.184U  W=8.026U
M6      U9_drain U8_drain VDD     VDD     P   L=0.18U  W=0.42U
M7      U8_drain U8_gate VSS     VSS     N   L=0.69U  W=0.24U
M8      U8_gate U6_gate VSS     VSS     N   L=1.16U  W=0.24U
M9      U1_drain I       VSS     VSS     N   L=0.18U  W=0.42U
M10     U6_gate U1_drain VSS     VSS     N   L=0.5U  W=0.24U
M11     U9_drain U8_drain VSS     VSS     N   L=0.18U  W=0.44U
M12     Z       U9_drain VSS     VSS     N   L=0.187U  W=3.30U

.ENDS dl03d4

.SUBCKT dl04d2 Z  I VDD VSS
M1      U8_drain U8_gate VDD     VDD     P   L=1.47U      W=0.42U
M2      U8_gate U6_gate VDD      VDD     P   L=2.76U      W=0.42U
M3      U1_drain I       VDD     VDD     P   L=0.18U      W=1.94U
M4      U6_gate U1_drain VDD     VDD     P   L=1.12U      W=0.42U
M5      Z       U9_drain VDD     VDD     P   L=0.187U     W=3.88U
M6      U9_drain U8_drain VDD    VDD     P   L=0.18U      W=0.42U
M7      U8_drain U8_gate VSS     VSS     N   L=1.25U      W=0.24U
M8      U8_gate U6_gate VSS      VSS     N   L=2.15U      W=0.24U
M9      U1_drain I       VSS     VSS     N   L=0.18U      W=0.42U
M10     U6_gate U1_drain VSS     VSS     N   L=0.76U      W=0.24U
M11     U9_drain U8_drain VSS    VSS     N   L=0.18U      W=0.37U
M12     Z       U9_drain VSS     VSS     N   L=0.18U      W=1.66U

.ENDS dl04d2

.SUBCKT dl04d4 Z  I VDD VSS
M1      U8_drain U8_gate VDD     VDD     P   L=1.47U  W=0.42U  
M2      U8_gate U6_gate VDD     VDD     P   L=2.75U  W=0.42U  
M3      U1_drain I       VDD     VDD     P   L=0.184U  W=1.94U  
M4      U6_gate U1_drain VDD     VDD     P   L=1.11U  W=0.42U  
M5      Z       U9_drain VDD     VDD     P   L=0.184U  W=8.2U  
M6      U9_drain U8_drain VDD     VDD     P   L=0.18U  W=0.42U  
M7      U8_drain U8_gate VSS     VSS     N   L=1.18U  W=0.24U  
M8      U8_gate U6_gate VSS     VSS     N   L=2.29U  W=0.24U  
M9      U1_drain I       VSS     VSS     N   L=0.18U  W=0.42U  
M10     U6_gate U1_drain VSS     VSS     N   L=0.76U  W=0.24U  
M11     U9_drain U8_drain VSS     VSS     N   L=0.18U  W=0.37U  
M12     Z       U9_drain VSS     VSS     N   L=0.18U  W=2.78U  

.ENDS dl04d4

.SUBCKT gclfsn1 GCLK  CLK EN SE VDD VSS
M1      u9_S    u9_GB   u9_D    VDD     P   L=0.18U    W=1.73U
M2      u9_S    u9_G    u9_D    VSS     N   L=0.18U      W=0.62U
M3      u9_D    u9_G    U23_out VDD     P   L=0.184U    W=1.73U
M4      u9_D    u9_GB   U23_out VSS     N   L=0.18U    W=0.62U
M5      GCLK    U34_in2 VDD     VDD     P   L=0.18U     W=2.08U
M6      GCLK    u9_G    VDD     VDD     P   L=0.184U    W=2.08U
M7      U34_$$7 U34_in2 VSS     VSS     N   L=0.18U     W=1.19U
M8      GCLK    u9_G    U34_$$7 VSS     N   L=0.18U     W=1.19U
M9      U34_in2 U32_out VDD     VDD     P   L=0.187U     W=1.50U
M10     U34_in2 u9_D    VDD     VDD     P   L=0.185U      W=1.50U
M11     U33_$$7 U32_out VSS     VSS     N   L=0.18U    W=0.84U
M12     U34_in2 u9_D    U33_$$7 VSS     N   L=0.18U      W=0.84U
M13     u9_S    U27_in  VSS     VSS     N   L=0.18U     W=0.62U
M14     u9_S    U27_in  VDD     VDD     P   L=0.184U    W=1.73U
M15     U27_in  u9_D    VSS     VSS     N   L=0.18U     W=0.62U
M16     U27_in  u9_D    VDD     VDD     P   L=0.184U     W=1.73U
M17     u9_GB   u9_G    VSS     VSS     N   L=0.18U    W=0.69U
M18     u9_GB   u9_G    VDD     VDD     P   L=0.184U    W=2.01U
M19     u9_G    CLK     VSS     VSS     N   L=0.18U     W=0.55U
M20     u9_G    CLK     VDD     VDD     P   L=0.184U    W=2.01U
M21     U23_out EN      VSS     VSS     N   L=0.18U     W=0.53U
M22     U23_out EN      VDD     VDD     P   L=0.18U      W=1.50U
M23     U32_out SE      VSS     VSS     N   L=0.18U     W=0.69U
M24     U32_out SE      VDD     VDD     P   L=0.184U     W=1.95U

.ENDS gclfsn1

.SUBCKT gclfsn2 GCLK  CLK EN SE VDD VSS
M1      u9_S    u9_GB   u9_D    VDD     P   L=0.184U  W=1.91U
M2      u9_S    u9_G    u9_D    VSS     N   L=0.18U   W=0.55U
M3      u9_D    u9_G    U23_out VDD     P   L=0.18U   W=1.86U
M4      u9_D    u9_GB   U23_out VSS     N   L=0.18U   W=0.62U
M5      u9_S    U27_in  VSS     VSS     N   L=0.18U   W=0.55U
M6      u9_S    U27_in  VDD     VDD     P   L=0.18U   W=1.73U
M7      u9_GB   u9_G    VSS     VSS     N   L=0.18U   W=0.83U
M8      u9_GB   u9_G    VDD     VDD     P   L=0.185U  W=1.83U
M9      u9_G    CLK     VSS     VSS     N   L=0.18U   W=0.62U    
M10     u9_G    CLK     VDD     VDD     P   L=0.184U  W=2.06U    
M11     U23_out EN      VSS     VSS     N   L=0.18U   W=0.42U  
M12     U23_out EN      VDD     VDD     P   L=0.185U  W=1.47U   
M13     U27_in  u9_D    VSS     VSS     N   L=0.18U   W=0.58U  
M14     U27_in  u9_D    VDD     VDD     P   L=0.184U  W=1.73U   
M15     GCLK    U30_out VSS     VSS     N   L=0.185U  W=1.5U  
M16     GCLK    U30_out VDD     VDD     P   L=0.1835U W=4.1U  
M17     U29_out SE      VSS     VSS     N   L=0.18U   W=0.42U   
M18     U29_out U27_in  VSS     VSS     N   L=0.18U   W=0.42U    
M19     U29_out U27_in  U29_$$7 VDD     P   L=0.183U  W=1.98U    
M20     U29_$$7 SE      VDD     VDD     P   L=0.183U  W=1.98U   
M21     U30_out U29_out VSS     VSS     N   L=0.18U   W=0.44U    
M22     U30_out u9_GB   VSS     VSS     N   L=0.18U   W=0.44U   
M23     U30_out u9_GB   U30_$$7 VDD     P   L=0.183U  W=2.33U   
M24     U30_$$7 U29_out VDD     VDD     P   L=0.183U  W=2.33U   

.ENDS gclfsn2

.SUBCKT gclfsn4 GCLK  CLK EN SE VDD VSS
M1      u9_S    u9_GB   u9_D    VDD     P   L=0.184U  W=1.91U  
M2      u9_S    u9_G    u9_D    VSS     N   L=0.18U  W=0.55U  
M3      u9_D    u9_G    U23_out VDD     P   L=0.18U  W=1.86U  
M4      u9_D    u9_GB   U23_out VSS     N   L=0.18U  W=0.62U  
M5      u9_S    U27_in  VSS     VSS     N   L=0.18U  W=0.55U  
M6      u9_S    U27_in  VDD     VDD     P   L=0.18U  W=1.73U  
M7      u9_GB   u9_G    VSS     VSS     N   L=0.18U  W=0.83U  
M8      u9_GB   u9_G    VDD     VDD     P   L=0.184U  W=1.83U  
M9      u9_G    CLK     VSS     VSS     N   L=0.18U  W=0.62U  
M10     u9_G    CLK     VDD     VDD     P   L=0.186U  W=2.1U  
M11     U23_out EN      VSS     VSS     N   L=0.18U  W=0.42U  
M12     U23_out EN      VDD     VDD     P   L=0.185U  W=1.47U  
M13     U27_in  u9_D    VSS     VSS     N   L=0.18U  W=0.58U  
M14     U27_in  u9_D    VDD     VDD     P   L=0.184U  W=1.73U  
M15     GCLK    U30_out VSS     VSS     N   L=0.18U  W=3.02U  
M16     GCLK    U30_out VDD     VDD     P   L=0.186U  W=7.09U  
M17     U29_out SE      VSS     VSS     N   L=0.18U  W=0.42U  
M18     U29_out U27_in  VSS     VSS     N   L=0.18U  W=0.42U  
M19     U29_out U27_in  U29_$$7 VDD     P   L=0.184U  W=1.98U  
M20     U29_$$7 SE      VDD     VDD     P   L=0.184U  W=1.98U  
M21     U30_out U29_out VSS     VSS     N   L=0.18U  W=0.44U  
M22     U30_out u9_GB   VSS     VSS     N   L=0.18U  W=0.44U  
M23     U30_out u9_GB   U30_$$7 VDD     P   L=0.183U  W=2.41U  
M24     U30_$$7 U29_out VDD     VDD     P   L=0.183U  W=2.41U  

.ENDS gclfsn4

.SUBCKT gclfsn7 GCLK  CLK EN SE VDD VSS
M1      u9_S    u9_GB   u9_D    VDD     P   L=0.184U  W=1.91U  
M2      u9_S    u9_G    u9_D    VSS     N   L=0.18U  W=0.55U  
M3      u9_D    u9_G    U23_out VDD     P   L=0.18U  W=1.86U  
M4      u9_D    u9_GB   U23_out VSS     N   L=0.18U  W=0.62U  
M5      u9_S    U27_in  VSS     VSS     N   L=0.18U  W=0.55U  
M6      u9_S    U27_in  VDD     VDD     P   L=0.18U  W=1.73U  
M7      u9_GB   u9_G    VSS     VSS     N   L=0.18U  W=0.83U  
M8      u9_GB   u9_G    VDD     VDD     P   L=0.184U  W=1.83U  
M9      u9_G    CLK     VSS     VSS     N   L=0.18U  W=0.62U  
M10     u9_G    CLK     VDD     VDD     P   L=0.186U  W=2.1U  
M11     U23_out EN      VSS     VSS     N   L=0.18U  W=0.42U  
M12     U23_out EN      VDD     VDD     P   L=0.185U  W=1.47U  
M13     U27_in  u9_D    VSS     VSS     N   L=0.18U  W=0.58U  
M14     U27_in  u9_D    VDD     VDD     P   L=0.184U  W=1.73U  
M15     GCLK    U30_out VSS     VSS     N   L=0.184U  W=5.23U  
M16     GCLK    U30_out VDD     VDD     P   L=0.182U  W=13.51U  
M17     U29_out SE      VSS     VSS     N   L=0.18U  W=0.42U  
M18     U29_out U27_in  VSS     VSS     N   L=0.18U  W=0.42U  
M19     U29_out U27_in  U29_$$7 VDD     P   L=0.184U  W=1.98U  
M20     U29_$$7 SE      VDD     VDD     P   L=0.184U  W=1.98U  
M21     U30_out U29_out VSS     VSS     N   L=0.18U  W=0.44U  
M22     U30_out u9_GB   VSS     VSS     N   L=0.18U  W=0.44U  
M23     U30_out u9_GB   U30_$$7 VDD     P   L=0.183U  W=2.51U  
M24     U30_$$7 U29_out VDD     VDD     P   L=0.183U  W=2.51U  

.ENDS gclfsn7

.SUBCKT gclfsna GCLK  CLK EN SE VDD VSS
M1      u9_S    u9_GB   u9_D    VDD     P   L=0.184U     W=1.91U
M2      u9_S    u9_G    u9_D    VSS     N   L=0.18U      W=0.55U
M3      u9_D    u9_G    U23_out VDD     P   L=0.18U      W=1.86U
M4      u9_D    u9_GB   U23_out VSS     N   L=0.18U      W=0.62U
M5      u9_S    U27_in  VSS     VSS     N   L=0.18U      W=0.55U
M6      u9_S    U27_in  VDD     VDD     P   L=0.18U      W=1.73U
M7      u9_GB   u9_G    VSS     VSS     N   L=0.18U      W=0.83U
M8      u9_GB   u9_G    VDD     VDD     P   L=0.184U     W=1.86U
M9      u9_G    CLK     VSS     VSS     N   L=0.18U      W=0.62U
M10     u9_G    CLK     VDD     VDD     P   L=0.184U     W=2.06U
M11     U23_out EN      VSS     VSS     N   L=0.18U      W=0.42U
M12     U23_out EN      VDD     VDD     P   L=0.185U     W=1.47U
M13     U27_in  u9_D    VSS     VSS     N   L=0.18U      W=0.58U
M14     U27_in  u9_D    VDD     VDD     P   L=0.184U     W=1.73U
M15     GCLK    U30_out VSS     VSS     N   L=0.18U     W=7.78U
M16     GCLK    U30_out VDD     VDD     P   L=0.18U      W=19.7U
M17     U29_out SE      VSS     VSS     N   L=0.18U      W=0.42U
M18     U29_out U27_in  VSS     VSS     N   L=0.18U      W=0.42U
M19     U29_out U27_in  U29_$$7 VDD     P   L=0.184U     W=1.98U
M20     U29_$$7 SE      VDD     VDD     P   L=0.184U     W=1.98U
M21     U30_out U29_out VSS     VSS     N   L=0.18U      W=0.83U
M22     U30_out u9_GB   VSS     VSS     N   L=0.18U      W=0.83U
M23     U30_out u9_GB   U30_$$7 VDD     P   L=0.184U     W=4.15U
M24     U30_$$7 U29_out VDD     VDD     P   L=0.182U     W=4.15U

.ENDS gclfsna

.SUBCKT gclrsn1 GCLK  CLK EN SE VDD VSS
M1      U24_out U24_in  VSS     VSS     N   L=0.18U  W=0.62U  
M2      U24_out U24_in  VDD     VDD     P   L=0.184U  W=1.91U  
M3      u9_GB   CLK     VSS     VSS     N   L=0.18U  W=0.55U  
M4      u9_GB   CLK     VDD     VDD     P   L=0.184U  W=2.06U  
M5      u9_G    u9_GB   VSS     VSS     N   L=0.18U  W=0.68U  
M6      u9_G    u9_GB   VDD     VDD     P   L=0.184U  W=1.73U  
M7      U23_out EN      VSS     VSS     N   L=0.18U  W=0.47U  
M8      U23_out EN      VDD     VDD     P   L=0.185U  W=1.3U  
M9      U24_in  QN      VSS     VSS     N   L=0.18U  W=0.62U  
M10     U24_in  QN      VDD     VDD     P   L=0.184U  W=1.91U  
M11     QN      u9_GB   U24_out VDD     P   L=0.18U  W=1.8U  
M12     QN      u9_G    U24_out VSS     N   L=0.18U  W=0.62U  
M13     U23_out u9_G    QN      VDD     P   L=0.184U  W=1.742U  
M14     U23_out u9_GB   QN      VSS     N   L=0.18U  W=0.62U  
M15     GCLK    U27_in1 VSS     VSS     N   L=0.18U  W=0.76U  
M16     GCLK    u9_GB   VSS     VSS     N   L=0.18U  W=0.76U  
M17     GCLK    u9_GB   U27_$$7 VDD     P   L=0.182U  W=3.95U  
M18     U27_$$7 U27_in1 VDD     VDD     P   L=0.182U  W=3.95U  
M19     U27_in1 SE      VSS     VSS     N   L=0.18U  W=0.42U  
M20     U27_in1 U24_in  VSS     VSS     N   L=0.18U  W=0.42U  
M21     U27_in1 U24_in  U26_$$7 VDD     P   L=0.18U  W=1.91U  
M22     U26_$$7 SE      VDD     VDD     P   L=0.18U  W=1.91U  

.ENDS gclrsn1

.SUBCKT gclrsn2 GCLK  CLK EN SE VDD VSS
M1      U24_out U24_in  VSS     VSS     N   L=0.18U     W=0.69U
M2      U24_out U24_in  VDD     VDD     P   L=0.18U    W=1.91U
M3      U24_in  QN      VSS     VSS     N   L=0.18U    W=0.69U
M4      U24_in  QN      VDD     VDD     P   L=0.184U     W=1.91U
M5      u9_GB   CLK     VSS     VSS     N   L=0.18U    W=0.62U
M6      u9_GB   CLK     VDD     VDD     P   L=0.184U     W=2.08U
M7      u9_G    u9_GB   VSS     VSS     N   L=0.18U    W=0.69U
M8      u9_G    u9_GB   VDD     VDD     P   L=0.184U     W=2.08U
M9      U23_out EN      VSS     VSS     N   L=0.18U     W=0.42U
M10     U23_out EN      VDD     VDD     P   L=0.185U     W=1.30U
M11     GCLK    U30_out VSS     VSS     N   L=0.185U    W=1.55U
M12     GCLK    U30_out VDD     VDD     P   L=0.182U      W=4.18U
M13     U28_out SE      VSS     VSS     N   L=0.18U     W=0.69U
M14     U28_out SE      VDD     VDD     P   L=0.184U     W=1.91U
M15     QN      u9_GB   U24_out VDD     P   L=0.184U     W=1.8U
M16     QN      u9_G    U24_out VSS     N   L=0.18U     W=0.62U
M17     U23_out u9_G    QN      VDD     P   L=0.18U     W=1.8U
M18     U23_out u9_GB   QN      VSS     N   L=0.18U    W=0.62U
M19     U30_out U30_in2 VDD     VDD     P   L=0.184U     W=1.87U
M20     U30_out u9_G    VDD     VDD     P   L=0.18U      W=1.87U
M21     U30_$$7 U30_in2 VSS     VSS     N   L=0.18U      W=0.97U
M22     U30_out u9_G    U30_$$7 VSS     N   L=0.18U     W=0.97U
M23     U30_in2 U28_out VDD     VDD     P   L=0.18U    W=1.91U
M24     U30_in2 QN      VDD     VDD     P   L=0.184U      W=1.91U
M25     U29_$$7 U28_out VSS     VSS     N   L=0.18U   W=0.69U
M26     U30_in2 QN      U29_$$7 VSS     N   L=0.18U    W=0.69U

.ENDS gclrsn2

.SUBCKT gclrsn4 GCLK  CLK EN SE VDD VSS
M1      U24_out U24_in  VSS     VSS     N   L=0.18U    W=0.69U
M2      U24_out U24_in  VDD     VDD     P   L=0.18U   W=1.91U
M3      U24_in  QN      VSS     VSS     N   L=0.18U     W=0.69U
M4      U24_in  QN      VDD     VDD     P   L=0.184U    W=1.91U
M5      u9_GB   CLK     VSS     VSS     N   L=0.18U     W=0.69U
M6      u9_GB   CLK     VDD     VDD     P   L=0.185U     W=2.08U
M7      u9_G    u9_GB   VSS     VSS     N   L=0.18U    W=0.69U
M8      u9_G    u9_GB   VDD     VDD     P   L=0.185U      W=2.08U
M9      U23_out EN      VSS     VSS     N   L=0.18U    W=0.42U
M10     U23_out EN      VDD     VDD     P   L=0.185U     W=1.30U
M11     GCLK    U30_out VSS     VSS     N   L=0.185U     W=3.32U
M12     GCLK    U30_out VDD     VDD     P   L=0.18U      W=8.64U
M13     U28_out SE      VSS     VSS     N   L=0.18U     W=0.69U
M14     U28_out SE      VDD     VDD     P   L=0.184U     W=1.91U
M15     QN      u9_GB   U24_out VDD     P   L=0.184U     W=1.8U
M16     QN      u9_G    U24_out VSS     N   L=0.18U      W=0.62U
M17     U23_out u9_G    QN      VDD     P   L=0.18U    W=1.8U
M18     U23_out u9_GB   QN      VSS     N   L=0.18U     W=0.62U
M19     U30_out U30_in2 VDD     VDD     P   L=0.184U    W=1.99U
M20     U30_out u9_G    VDD     VDD     P   L=0.18U     W=1.99U
M21     U30_$$7 U30_in2 VSS     VSS     N   L=0.18U     W=1U
M22     U30_out u9_G    U30_$$7 VSS     N   L=0.18U     W=1U
M23     U30_in2 U28_out VDD     VDD     P   L=0.18U     W=1.91U
M24     U30_in2 QN      VDD     VDD     P   L=0.184U      W=1.91U
M25     U29_$$7 U28_out VSS     VSS     N   L=0.18U     W=0.69U
M26     U30_in2 QN      U29_$$7 VSS     N   L=0.18U    W=0.69U

.ENDS gclrsn4

.SUBCKT gclrsn7 GCLK  CLK EN SE VDD VSS
M1      U24_out U24_in  VSS     VSS     N   L=0.18U     W=0.69U
M2      U24_out U24_in  VDD     VDD     P   L=0.18U    W=1.91U
M3      U24_in  QN      VSS     VSS     N   L=0.18U      W=0.69U
M4      U24_in  QN      VDD     VDD     P   L=0.184U      W=1.91U
M5      u9_GB   CLK     VSS     VSS     N   L=0.18U      W=0.692U
M6      u9_GB   CLK     VDD     VDD     P   L=0.184U      W=2.08U
M7      u9_G    u9_GB   VSS     VSS     N   L=0.18U      W=0.69U
M8      u9_G    u9_GB   VDD     VDD     P   L=0.184U      W=2.08U
M9      U23_out EN      VSS     VSS     N   L=0.18U    W=0.42U
M10     U23_out EN      VDD     VDD     P   L=0.186U     W=1.30U
M11     GCLK    U30_out VSS     VSS     N   L=0.184U     W=5.54U
M12     GCLK    U30_out VDD     VDD     P   L=0.18U     W=13.42U
M13     U28_out SE      VSS     VSS     N   L=0.18U      W=0.69U
M14     U28_out SE      VDD     VDD     P   L=0.184U     W=1.91U
M15     QN      u9_GB   U24_out VDD     P   L=0.184U     W=1.8U
M16     QN      u9_G    U24_out VSS     N   L=0.18U     W=0.6223U
M17     U23_out u9_G    QN      VDD     P   L=0.18U      W=1.8U
M18     U23_out u9_GB   QN      VSS     N   L=0.18U     W=0.62U
M19     U30_out U30_in2 VDD     VDD     P   L=0.184U      W=2.13U
M20     U30_out u9_G    VDD     VDD     P   L=0.18U      W=2.13U
M21     U30_$$7 U30_in2 VSS     VSS     N   L=0.18U     W=1.11U
M22     U30_out u9_G    U30_$$7 VSS     N   L=0.18U    W=1.11U
M23     U30_in2 U28_out VDD     VDD     P   L=0.18U     W=1.91U
M24     U30_in2 QN      VDD     VDD     P   L=0.184U      W=1.91U
M25     U29_$$7 U28_out VSS     VSS     N   L=0.18U      W=0.69U
M26     U30_in2 QN      U29_$$7 VSS     N   L=0.18U     W=0.69U

.ENDS gclrsn7

.SUBCKT gclrsna GCLK  CLK EN SE VDD VSS
M1      U24_out U24_in  VSS     VSS     N   L=0.18U     W=0.69U
M2      U24_out U24_in  VDD     VDD     P   L=0.18U     W=1.91U
M3      U24_in  QN      VSS     VSS     N   L=0.18U    W=0.69U
M4      U24_in  QN      VDD     VDD     P   L=0.184U    W=1.91U
M5      u9_GB   CLK     VSS     VSS     N   L=0.18U    W=0.69U
M6      u9_GB   CLK     VDD     VDD     P   L=0.184U    W=2.08U
M7      u9_G    u9_GB   VSS     VSS     N   L=0.18U   W=0.69U
M8      u9_G    u9_GB   VDD     VDD     P   L=0.184U  W=2.08U
M9      u8_S    EN      VSS     VSS     N   L=0.18U      W=0.42U
M10     u8_S    EN      VDD     VDD     P   L=0.186U    W=1.30U
M11     GCLK    U30_out VSS     VSS     N   L=0.187U     W=7.08U
M12     GCLK    U30_out VDD     VDD     P   L=0.182U      W=19.09U
M13     U28_out SE      VSS     VSS     N   L=0.18U     W=0.69U
M14     U28_out SE      VDD     VDD     P   L=0.184U     W=1.91U
M15     QN      u9_GB   U24_out VDD     P   L=0.184U      W=1.8U
M16     QN      u9_G    U24_out VSS     N   L=0.18U      W=0.62U
M17     u8_S    u9_G    QN      VDD     P   L=0.18U      W=1.8U
M18     u8_S    u9_GB   QN      VSS     N   L=0.18U      W=0.62U
M19     U30_out U30_in2 VDD     VDD     P   L=0.184U      W=2.13U
M20     U30_out u9_G    VDD     VDD     P   L=0.18U      W=2.13U
M21     U30_$$7 U30_in2 VSS     VSS     N   L=0.18U      W=1.22U
M22     U30_out u9_G    U30_$$7 VSS     N   L=0.18U      W=1.22U
M23     U30_in2 U28_out VDD     VDD     P   L=0.18U      W=1.91U
M24     U30_in2 QN      VDD     VDD     P   L=0.184U      W=1.91U
M25     U29_$$7 U28_out VSS     VSS     N   L=0.18U      W=0.69U
M26     U30_in2 QN      U29_$$7 VSS     N   L=0.18U      W=0.69U

.ENDS gclrsna

.SUBCKT gcnfnn1 GCLK  CLK EN VDD VSS
M1      U3_drain EN      VDD     VDD     P   L=0.184U  W=1.65U   
+  PD=.820U
M2      U3_drain CLK     VDD     VDD     P   L=0.185U  W=1.62U   
+  PD=.820U
M3      GCLK    U3_drain VDD     VDD     P   L=0.184U  W=2.06U   
+  PD=1.505U
M4      u2_drain EN      VSS     VSS     N   L=0.18U  W=0.66U   
+  PD=.700U
M5      U3_drain CLK     u2_drain VSS     N   L=0.18U  W=0.66U   
+  PS=.700U PD=.700U
M6      GCLK    U3_drain VSS     VSS     N   L=0.18U  W=0.75U   
+  PD=1.382U

.ENDS gcnfnn1

.SUBCKT gcnfnn2 GCLK  CLK EN VDD VSS
M1      U3_drain EN      VDD     VDD     P   L=0.185U  W=1.69U   
+  PD=.820U
M2      U3_drain CLK     VDD     VDD     P   L=0.185U  W=1.63U   
+  PD=.820U
M3      GCLK    U3_drain VDD     VDD     P   L=0.1845U  W=4.38U   
+  PD=1.505U
M4      u2_drain EN      VSS     VSS     N   L=0.18U  W=0.66U   
+  PD=.700U
M5      U3_drain CLK     u2_drain VSS     N   L=0.18U  W=0.66U   
+  PS=.700U PD=.700U
M6      GCLK    U3_drain VSS     VSS     N   L=0.186U  W=1.36U   
+  PD=1.382U

.ENDS gcnfnn2

.SUBCKT gcnfnn4 GCLK  CLK EN VDD VSS
M1      U3_drain EN      VDD     VDD     P   L=0.18U       W=2.22U
+  PD=.820U
M2      U3_drain CLK     VDD     VDD     P   L=0.186U      W=2.102U
+  PD=.820U
M3      GCLK    U3_drain VDD     VDD     P   L=0.18U       W=8.86U
+  PD=1.505U
M4      u2_drain EN      VSS     VSS     N   L=0.18U       W=0.9U
+  PD=.700U
M5      U3_drain CLK     u2_drain VSS     N   L=0.18U      W=0.9U
+  PS=.700U PD=.700U
M6      GCLK    U3_drain VSS     VSS     N   L=0.18U       W=2.99U
+  PD=1.382U

.ENDS gcnfnn4

.SUBCKT gcnfnn7 GCLK  CLK EN VDD VSS
M1      U3_drain EN      VDD     VDD     P   L=0.184U  W=2.07U   
+  PD=.820U
M2      U3_drain CLK     VDD     VDD     P   L=0.18U  W=2.33U   
+  PD=.820U
M3      GCLK    U3_drain VDD     VDD     P   L=0.185167U  W=14.34U   
+  PD=1.505U
M4      u2_drain EN      VSS     VSS     N   L=0.18U  W=1U   
+  PD=.700U
M5      U3_drain CLK     u2_drain VSS     N   L=0.18U  W=1U   
+  PS=.700U PD=.700U
M6      GCLK    U3_drain VSS     VSS     N   L=0.1824U  W=5.12U   
+  PD=1.382U

.ENDS gcnfnn7

.SUBCKT gcnfnna GCLK  CLK EN VDD VSS
M1      U3_drain EN      VDD     VDD     P   L=0.18U       W=2.26U
+  PD=.820U
M2      U3_drain CLK     VDD     VDD     P   L=0.184U       W=2.069U
+  PD=.820U
M3      GCLK    U3_drain VDD     VDD     P   L=0.182U       W=19.88U
+  PD=1.505U
M4      u2_drain EN      VSS     VSS     N   L=0.18U       W=1.02U
+  PD=.700U
M5      U3_drain CLK     u2_drain VSS     N   L=0.18U       W=1.02U
+  PS=.700U PD=.700U
M6      GCLK    U3_drain VSS     VSS     N   L=0.18U       W=7.31U
+  PD=1.382U

.ENDS gcnfnna

.SUBCKT gcnrnn1 GCLK  CLK EN VDD VSS
M1      u2_drain EN      VSS     VSS     N   L=0.186U  W=1.34U   
+  PD=.700U
M2      GCLK    U4_gate u2_drain VSS     N   L=0.186U  W=1.34U   
+  PS=.700U PD=.700U
M3      GCLK    U4_gate VDD     VDD     P   L=0.183U  W=2.13U   PD=.820U
M4      GCLK    EN      VDD     VDD     P   L=0.183U  W=2.13U   PD=.820U
M5      U4_gate CLK     VSS     VSS     N   L=0.18U  W=0.55U  
M6      U4_gate CLK     VDD     VDD     P   L=0.184U  W=1.94U  

.ENDS gcnrnn1

.SUBCKT gcnrnn2 GCLK  CLK EN VDD VSS
M1      GCLK    U39_in  VSS     VSS     N   L=0.18U  W=1.77U  
M2      GCLK    U39_in  VDD     VDD     P   L=0.1835U  W=4.85U  
M3      u2_gate EN      VSS     VSS     N   L=0.18U  W=0.44U  
M4      u2_gate EN      VDD     VDD     P   L=0.186U  W=1.30U  
M5      U39_in  u2_gate VSS     VSS     N   L=0.18U  W=0.44U   PD=.430U
M6      U39_in  CLK     VSS     VSS     N   L=0.18U  W=0.44U   PD=.430U
M7      U39_in  CLK     u1_source VDD     P   L=0.183U  W=2.59U   
+  PS=.840U PD=.840U
M8      VDD     u2_gate u1_source VDD     P   L=0.183U  W=2.59U   
+  PS=.840U

.ENDS gcnrnn2

.SUBCKT gcnrnn4 GCLK  CLK EN VDD VSS
M1      GCLK    U39_in  VSS     VSS     N   L=0.18U  W=3.16U  
M2      GCLK    U39_in  VDD     VDD     P   L=0.182U  W=8.72U  
M3      u2_gate EN      VSS     VSS     N   L=0.18U  W=0.50U  
M4      u2_gate EN      VDD     VDD     P   L=0.184U  W=2.01U  
M5      U39_in  u2_gate VSS     VSS     N   L=0.18U  W=0.42U   PD=.430U
M6      U39_in  CLK     VSS     VSS     N   L=0.18U  W=0.42U   PD=.430U
M7      U39_in  CLK     u1_source VDD     P   L=0.18U  W=2.63U   
+  PS=.840U PD=.840U
M8      VDD     u2_gate u1_source VDD     P   L=0.18U  W=2.63U   
+  PS=.840U

.ENDS gcnrnn4

.SUBCKT gcnrnn7 GCLK  CLK EN VDD VSS
M1      GCLK    U39_in  VSS     VSS     N   L=0.18U  W=5.23U  
M2      GCLK    U39_in  VDD     VDD     P   L=0.18U  W=12.67U  
M3      u2_gate EN      VSS     VSS     N   L=0.18U  W=0.62U  
M4      u2_gate EN      VDD     VDD     P   L=0.184U  W=2.01U  
M5      U39_in  u2_gate VSS     VSS     N   L=0.18U  W=0.44U   PD=.430U
M6      U39_in  CLK     VSS     VSS     N   L=0.18U  W=0.44U   PD=.430U
M7      U39_in  CLK     u1_source VDD     P   L=0.183U  W=2.55U   
+  PS=.840U PD=.840U
M8      VDD     u2_gate u1_source VDD     P   L=0.183U  W=2.55U   
+  PS=.840U

.ENDS gcnrnn7

.SUBCKT gcnrnna GCLK  CLK EN VDD VSS
M1      GCLK    U39_in  VSS     VSS     N   L=0.18U  W=8.10U  
M2      GCLK    U39_in  VDD     VDD     P   L=0.182444U  W=20.28U  
M3      u2_gate EN      VSS     VSS     N   L=0.18U  W=0.62U  
M4      u2_gate EN      VDD     VDD     P   L=0.184U  W=2.01U  
M5      U39_in  u2_gate VSS     VSS     N   L=0.18U  W=0.44U   PD=.430U
M6      U39_in  CLK     VSS     VSS     N   L=0.18U  W=0.44U   PD=.430U
M7      U39_in  CLK     u1_source VDD     P   L=0.18U  W=2.58U   
+  PS=.840U PD=.840U
M8      VDD     u2_gate u1_source VDD     P   L=0.18U  W=2.58U   
+  PS=.840U

.ENDS gcnrnna

.SUBCKT invbd7 ZN  I VDD VSS
M1      ZN      I       VSS     VSS     N   L=0.180U    W=5.32U
M2      ZN      I       VDD     VDD     P   L=0.183U      W=14.82U

.ENDS invbd7

.SUBCKT invbda ZN  I VDD VSS
M1      ZN      I       VSS     VSS     N   L=0.18U      W=6.98U
M2      ZN      I       VDD     VDD     P   L=0.182333U   W=20.13U

.ENDS invbda

.SUBCKT invbdf ZN  I VDD VSS
M1      ZN      I       VSS     VSS     N   L=0.184455U  W=10.63U  
M2      ZN      I       VDD     VDD     P   L=0.183U  W=29.68U  

.ENDS invbdf

.SUBCKT invbdk ZN  I VDD VSS
M1      ZN      I       VSS     VSS     N   L=0.184U  W=14.18U  
M2      ZN      I       VDD     VDD     P   L=0.183938U  W=40.69U  

.ENDS invbdk

.SUBCKT jkbrb4 Q QN  CDN CP J KZ SDN VDD VSS
M1      U80_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.78U
M2      U80_out U80_in1 U80_u7_drain VSS     N   L=0.18U  W=0.78U
M3      U80_out U80_in1 VDD     VDD     P   L=0.18U  W=1.18U
M4      VDD     CDN     U80_out VDD     P   L=0.187U  W=1.18U
M5      U24_u7_drain U24_in2 VSS     VSS     N   L=0.18U  W=0.78U
M6      U80_in1 SDN     U24_u7_drain VSS     N   L=0.18U  W=0.78U
M7      U80_in1 SDN     VDD     VDD     P   L=0.187U  W=1.18U
M8      VDD     U24_in2 U80_in1 VDD     P   L=0.18U  W=1.18U
M9      U82_u7_drain U21_in  VSS     VSS     N   L=0.18U  W=0.78U
M10     U77_gate SDN     U82_u7_drain VSS     N   L=0.18U  W=0.78U
M11     U77_gate SDN     VDD     VDD     P   L=0.187U  W=1.11U
M12     VDD     U21_in  U77_gate VDD     P   L=0.187U  W=1.11U
M13     U81_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.78U
M14     U21_in  u8_D    U81_u7_drain VSS     N   L=0.18U  W=0.78U
M15     U21_in  u8_D    VDD     VDD     P   L=0.18U  W=0.99U
M16     VDD     CDN     U21_in  VDD     P   L=0.187U  W=1.11U
M17     U80_in1 u8_GB   u8_D    VDD     P   L=0.18U  W=1.08U
M18     U80_in1 u8_G    u8_D    VSS     N   L=0.18U  W=0.42U
M19     U15_S   u8_G    U24_in2 VDD     P   L=0.18U W=1.43U
M20     U15_S   u8_GB   U24_in2 VSS     N   L=0.18U  W=0.5U
M21     U80_out u8_GB   U24_in2 VDD     P   L=0.186U  W=1.29U
M22     U80_out u8_G    U24_in2 VSS     N   L=0.18U  W=0.55U
M23     U77_gate u8_G    u8_D    VDD     P   L=0.18U  W=0.84U
M24     U77_gate u8_GB   u8_D    VSS     N   L=0.18U  W=0.42U
M25     U76_drain KZ      U15_S   VSS     N   L=0.18U  W=0.6U
M26     U76_drain J       VSS     VSS     N   L=0.18U  W=0.58U
M27     U76_drain U77_gate VSS     VSS     N   L=0.18U  W=0.6U
M28     U15_S   U75_gate U76_drain VSS     N   L=0.18U  W=0.58U
M29     Q       U21_in  VSS     VSS     N   L=0.18U  W=2.99U
M30     Q       U21_in  VDD     VDD     P   L=0.18375U  W=8.31U
M31     u8_GB   CP      VSS     VSS     N   L=0.18U  W=0.46U
M32     u8_GB   CP      VDD     VDD     P   L=0.18U  W=1.04U
M33     u8_G    u8_GB   VSS     VSS     N   L=0.18U  W=0.46U
M34     u8_G    u8_GB   VDD     VDD     P   L=0.18U  W=1.04U
M35     U75_gate U77_gate VSS     VSS     N   L=0.18U  W=0.58U
M36     U75_gate U77_gate VDD     VDD     P   L=0.185U  W=1.49U
M37     QN      u8_D    VSS     VSS     N   L=0.18U W=2.82U
M38     QN      u8_D    VDD     VDD     P   L=0.182U  W=8.31U
M39     U15_S   KZ      U73_source VDD     P   L=0.18U  W=1.44U
M40     U73_source U75_gate VDD     VDD     P   L=0.18U  W=1.44U
M41     u17_drain J       U15_S   VDD     P   L=0.18U  W=1.44U
M42     VDD     U77_gate u17_drain VDD     P   L=0.18U  W=1.44U

.ENDS jkbrb4

.SUBCKT labhb4 Q QN  CDN D E SDN VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.184U     W=1.77U
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U     W=0.69U
M3      u9_S    u8_G    u8_S    VDD     P   L=0.186U      W=1.77U
M4      u9_S    u8_GB   u8_S    VSS     N   L=0.18U      W=0.69U
M5      QN      U22_in  VSS     VSS     N   L=0.18U      W=2.91U
M6      QN      U22_in  VDD     VDD     P   L=0.18275U      W=8.2U
M7      u8_G    u8_GB   VSS     VSS     N   L=0.18U      W=0.69U
M8      u8_G    u8_GB   VDD     VDD     P   L=0.18U     W=1.77U
M9      u8_GB   E       VSS     VSS     N   L=0.18U      W=0.69U
M10     u8_GB   E       VDD     VDD     P   L=0.184U      W=1.77U
M11     U22_in  u9_S    VSS     VSS     N   L=0.18U      W=0.69U
M12     U22_in  u9_S    VDD     VDD     P   L=0.184U      W=2.05U
M13     u3_out  u3_in   VSS     VSS     N   L=0.18U      W=0.61U
M14     u3_out  u3_in   VDD     VDD     P   L=0.18U      W=1.56U
M15     Q       u3_out  VSS     VSS     N   L=0.18U      W=2.91U
M16     Q       u3_out  VDD     VDD     P   L=0.18U      W=8.2U
M17     U26_u7_drain D       VSS     VSS     N   L=0.18U      W=0.66U
M18     u8_D    CDN     U26_u7_drain VSS     N   L=0.18U      W=0.66U
M19     u8_D    CDN     VDD     VDD     P   L=0.18U      W=1.66U
M20     VDD     D       u8_D    VDD     P   L=0.185U      W=1.7U
M21     U24_u7_drain SDN     VSS     VSS     N   L=0.18U      W=1.11U
M22     u3_in   u8_S    U24_u7_drain VSS     N   L=0.18U      W=1.11U
M23     u3_in   u8_S    VDD     VDD     P   L=0.185U      W=1.7U
M24     VDD     SDN     u3_in   VDD     P   L=0.18U      W=1.7U
M25     U25_u7_drain u3_in   VSS     VSS     N   L=0.18U      W=1.11U
M26     u9_S    CDN     U25_u7_drain VSS     N   L=0.18U      W=1.11U
M27     u9_S    CDN     VDD     VDD     P   L=0.18U      W=1.65U
M28     VDD     u3_in   u9_S    VDD     P   L=0.185U      W=1.7U

.ENDS labhb4

.SUBCKT lachq4 Q  CDN D E VDD VSS
M1      u9_S         u9_GB   u9_D          VDD     P   L=0.184U  W=1.77U  
M2      u9_S         u9_G    u9_D          VSS     N   L=0.18U   W=0.73U  
M3      u9_D         u9_G    U29_out       VDD     P   L=0.183U  W=1.77U  
M4      u9_D         u9_GB   U29_out       VSS     N   L=0.18U   W=0.73U  
M5      u9_GB        u9_G    VSS           VSS     N   L=0.18U   W=0.69U  
M6      u9_GB        u9_G    VDD           VDD     P   L=0.184U  W=1.77U  
M7      u9_G         E       VSS           VSS     N   L=0.18U   W=0.69U  
M8      u9_G         E       VDD           VDD     P   L=0.184U  W=1.77U  
M9      Q            u9_D    VSS           VSS     N   L=0.18U   W=2.91U  
M10     Q            u9_D    VDD           VDD     P   L=0.183U  W=8.2U  
M11     U24_in2      u9_D    VSS           VSS     N   L=0.18U   W=0.77U  
M12     U24_in2      u9_D    VDD           VDD     P   L=0.185U  W=2.05U  
M13     U29_u7_drain D       VSS           VSS     N   L=0.18U   W=0.69U  
M14     U29_out      CDN     U29_u7_drain  VSS     N   L=0.18U   W=0.69U  
M15     U29_out      CDN     VDD           VDD     P   L=0.184U  W=1.72U  
M16     VDD          D       U29_out       VDD     P   L=0.184U  W=1.73U  
M17     U24_u7_drain U24_in2 VSS           VSS     N   L=0.18U   W=1.11U  
M18     u9_S         CDN     U24_u7_drain  VSS     N   L=0.18U   W=1.11U  
M19     u9_S         CDN     VDD           VDD     P   L=0.184U  W=1.65U  
M20     VDD          U24_in2 u9_S          VDD     P   L=0.184U  W=1.65U  

.ENDS lachq4

.SUBCKT laclq4 Q  CDN D EN VDD VSS
M1      u9_S    u9_GB   u9_D    VDD     P   L=0.184U  W=1.77U
M2      u9_S    u9_G    u9_D    VSS     N   L=0.18U  W=0.69U
M3      u8_S    u9_G    u9_S    VDD     P   L=0.184U  W=1.77U
M4      u8_S    u9_GB   u9_S    VSS     N   L=0.18U  W=0.69U
M5      U28_out u9_S    VSS     VSS     N   L=0.18U  W=0.77U
M6      U28_out u9_S    VDD     VDD     P   L=0.184U  W=2.05U
M7      u9_G    u9_GB   VSS     VSS     N   L=0.18U  W=0.69U
M8      u9_G    u9_GB   VDD     VDD     P   L=0.184U  W=1.73U
M9      u9_GB   EN      VSS     VSS     N   L=0.18U  W=0.69U
M10     u9_GB   EN      VDD     VDD     P   L=0.184U  W=1.73U
M11     Q       u9_S    VSS     VSS     N   L=0.18U  W=2.91U
M12     Q       u9_S    VDD     VDD     P   L=0.183U  W=8.2U
M13     U24_u7_drain D       VSS     VSS     N   L=0.18U  W=0.69U
M14     u8_S    CDN     U24_u7_drain VSS     N   L=0.18U  W=0.69U
M15     u8_S    CDN     VDD     VDD     P   L=0.184U  W=1.77U
M16     VDD     D       u8_S    VDD     P   L=0.184U  W=1.77U
M17     U29_u7_drain U28_out VSS     VSS     N   L=0.187U  W=1.11U
M18     u9_D    CDN     U29_u7_drain VSS     N   L=0.187U  W=1.11U
M19     u9_D    CDN     VDD     VDD     P   L=0.184U  W=1.74U
M20     VDD     U28_out u9_D    VDD     P   L=0.187U  W=1.7U

.ENDS laclq4

.SUBCKT lanhb4 Q QN  D E VDD VSS
M1      u9_S    u9_GB   u9_D    VDD     P   L=0.18U  W=1.08U  
M2      u9_S    u9_G    u9_D    VSS     N   L=0.18U  W=0.69U  
M3      u9_D    u9_G    u8_D    VDD     P   L=0.185U  W=1.73U  
M4      u9_D    u9_GB   u8_D    VSS     N   L=0.18U  W=0.42U  
M5      u9_GB   u9_G    VSS     VSS     N   L=0.18U  W=0.69U  
M6      u9_GB   u9_G    VDD     VDD     P   L=0.185U  W=1.715U  
M7      u9_G    E       VSS     VSS     N   L=0.18U  W=0.6U  
M8      u9_G    E       VDD     VDD     P   L=0.185U  W=1.47U  
M9      u8_D    D       VSS     VSS     N   L=0.18U  W=0.42U  
M10     u8_D    D       VDD     VDD     P   L=0.18U  W=1.08U  
M11     Q       u9_D    VSS     VSS     N   L=0.183U  W=2.88U  
M12     Q       u9_D    VDD     VDD     P   L=0.184U  W=8.18U  
M13     u9_S    U25_in  VSS     VSS     N   L=0.18U  W=0.69U  
M14     u9_S    U25_in  VDD     VDD     P   L=0.184U  W=1.77U  
M15     U25_in  u9_D    VSS     VSS     N   L=0.18U  W=0.69U  
M16     U25_in  u9_D    VDD     VDD     P   L=0.18U  W=1.77U  
M17     QN      U25_in  VSS     VSS     N   L=0.18U  W=2.88U  
M18     QN      U25_in  VDD     VDD     P   L=0.183667U  W=8.2U  

.ENDS lanhb4

.SUBCKT lanhn4 QN  D E VDD VSS
M1      u9_S    u9_GB   u9_D    VDD     P   L=0.186U  W=1.08U
M2      u9_S    u9_G    u9_D    VSS     N   L=0.18U  W=0.69U
M3      u9_D    u9_G    u8_D    VDD     P   L=0.185U  W=1.69U
M4      u9_D    u9_GB   u8_D    VSS     N   L=0.18U  W=0.42U
M5      u9_GB   u9_G    VSS     VSS     N   L=0.18U  W=0.69U
M6      u9_GB   u9_G    VDD     VDD     P   L=0.185U  W=1.66U
M7      u9_G    E       VSS     VSS     N   L=0.18U  W=0.5U
M8      u9_G    E       VDD     VDD     P   L=0.186U  W=1.29U
M9      U16_out D       VSS     VSS     N   L=0.18U  W=0.42U
M10     U16_out D       VDD     VDD     P   L=0.188U  W=1.04U
M11     u8_D    U16_out VSS     VSS     N   L=0.18U  W=0.42U
M12     u8_D    U16_out VDD     VDD     P   L=0.188U  W=1.04U
M13     QN      u9_D    VSS     VSS     N   L=0.1853U  W=2.91U
M14     QN      u9_D    VDD     VDD     P   L=0.183U  W=8.31U
M15     u9_S    U26_in  VSS     VSS     N   L=0.18U  W=0.69U
M16     u9_S    U26_in  VDD     VDD     P   L=0.18U  W=1.77U
M17     U26_in  u9_D    VSS     VSS     N   L=0.18U  W=0.69U
M18     U26_in  u9_D    VDD     VDD     P   L=0.184U  W=1.77U

.ENDS lanhn4

.SUBCKT lanhq4 Q  D E VDD VSS
M1      u9_S    u9_GB   u9_D    VDD     P   L=0.18U  W=1.08U  
M2      u9_S    u9_G    u9_D    VSS     N   L=0.18U  W=0.69U  
M3      u9_D    u9_G    U23_out VDD     P   L=0.184U  W=1.73U  
M4      u9_D    u9_GB   U23_out VSS     N   L=0.18U  W=0.42U  
M5      u9_GB   u9_G    VSS     VSS     N   L=0.18U  W=0.69U  
M6      u9_GB   u9_G    VDD     VDD     P   L=0.185U  W=1.73U  
M7      u9_G    E       VSS     VSS     N   L=0.18U  W=0.6U  
M8      u9_G    E       VDD     VDD     P   L=0.185U  W=1.43U  
M9      U23_out D       VSS     VSS     N   L=0.18U  W=0.42U  
M10     U23_out D       VDD     VDD     P   L=0.18U  W=1.08U  
M11     u9_S    U27_in  VSS     VSS     N   L=0.18U  W=0.69U  
M12     u9_S    U27_in  VDD     VDD     P   L=0.184U  W=1.77U  
M13     U27_in  u9_D    VSS     VSS     N   L=0.18U  W=0.69U  
M14     U27_in  u9_D    VDD     VDD     P   L=0.184U  W=1.77U  
M15     Q       u9_D    VSS     VSS     N   L=0.187U  W=2.91U  
M16     Q       u9_D    VDD     VDD     P   L=0.183U  W=8.24U  

.ENDS lanhq4

.SUBCKT lanht4 Z  D E OE VDD VSS
M1      U4_drain U4_gate U4_source VDD     P   L=0.18U       W=1.77U
+  PS=1.227U PD=1.145U
M2      U4_source U28_out VDD     VDD     P   L=0.184U       W=1.91U
+  PD=1.227U
M3      U4_source OE      VDD     VDD     P   L=0.18U       W=1.77U
+  PD=1.227U
M4      Z       U4_source VDD     VDD     P   L=0.1835U       W=4.1U
+  PD=2.018U
M5      Z       U4_source VDD     VDD     P   L=0.18U       W=4.1U
+  PD=2.018U
M6      U4_source OE      U4_drain VSS     N   L=0.18U       W=0.69U
+  PS=1.164U PD=1.239U
M7      Z       U4_drain VSS     VSS     N   L=0.18U       W=1.45U
+  PD=1.330U
M8      U4_drain U4_gate VSS     VSS     N   L=0.18U       W=0.69U
+  PD=1.164U
M9      U4_drain U28_out VSS     VSS     N   L=0.18U       W=0.69U
+  PD=1.164U
M10     Z       U4_drain VSS     VSS     N   L=0.18U       W=1.45U
+  PD=1.330U
M11     u11_out u11_in  VSS     VSS     N   L=0.18U      W=0.69U
M12     u11_out u11_in  VDD     VDD     P   L=0.185U      W=1.7U
M13     u11_in  E       VSS     VSS     N   L=0.18U      W=0.5U
M14     u11_in  E       VDD     VDD     P   L=0.18U      W=1.29U
M15     U4_gate OE      VSS     VSS     N   L=0.18U      W=0.69U
M16     U4_gate OE      VDD     VDD     P   L=0.18U      W=1.77U
M17     U28_out u8_S    VSS     VSS     N   L=0.18U      W=0.69U
M18     U28_out u8_S    VDD     VDD     P   L=0.18U      W=1.77U
M19     u8_D    D       VSS     VSS     N   L=0.18U      W=0.42U
M20     u8_D    D       VDD     VDD     P   L=0.18U      W=1.08U
M21     u9_S    U28_out VSS     VSS     N   L=0.18U      W=0.69U
M22     u9_S    U28_out VDD     VDD     P   L=0.185U      W=1.77U
M23     u8_S    u11_in  u8_D    VDD     P   L=0.184U      W=1.73U
M24     u8_S    u11_out u8_D    VSS     N   L=0.18U      W=0.42U
M25     u9_S    u11_out u8_S    VDD     P   L=0.18U      W=1.08U
M26     u9_S    u11_in  u8_S    VSS     N   L=0.18U      W=0.69U

.ENDS lanht4

.SUBCKT lanlb4 Q QN  D EN VDD VSS
M1      u9_S    u9_GB   u9_D    VDD     P   L=0.187U    W=1.08U  
M2      u9_S    u9_G    u9_D    VSS     N   L=0.18U     W=0.69U  
M3      u8_S    u9_G    u9_S    VDD     P   L=0.184U    W=1.77U  
M4      u8_S    u9_GB   u9_S    VSS     N   L=0.18U     W=0.42U  
M5      u9_G    u9_GB   VSS     VSS     N   L=0.18U     W=0.69U  
M6      u9_G    u9_GB   VDD     VDD     P   L=0.18U     W=1.73U  
M7      u9_GB   EN      VSS     VSS     N   L=0.18U     W=0.6U  
M8      u9_GB   EN      VDD     VDD     P   L=0.18U     W=1.43U  
M9      u8_S    D       VSS     VSS     N   L=0.18U     W=0.42U  
M10     u8_S    D       VDD     VDD     P   L=0.18U     W=1.08U  
M11     u9_D    U24_in  VSS     VSS     N   L=0.18U     W=0.69U  
M12     u9_D    U24_in  VDD     VDD     P   L=0.18U     W=1.77U  
M13     U24_in  u9_S    VSS     VSS     N   L=0.18U     W=0.69U  
M14     U24_in  u9_S    VDD     VDD     P   L=0.184U    W=1.78U  
M15     Q       u9_S    VSS     VSS     N   L=0.18U     W=2.94U  
M16     Q       u9_S    VDD     VDD     P   L=0.184U    W=8.18U  
M17     QN      U24_in  VSS     VSS     N   L=0.18U     W=2.94U  
M18     QN      U24_in  VDD     VDD     P   L=0.182U     W=8.2U  

.ENDS lanlb4

.SUBCKT lanln4 QN  D EN VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.185U  W=1.77U  
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U  W=0.42U  
M3      u8_D    u8_G    U26_out VDD     P   L=0.18U  W=1.04U  
M4      u8_D    u8_GB   U26_out VSS     N   L=0.18U  W=0.69U  
M5      u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.69U  
M6      u8_GB   u8_G    VDD     VDD     P   L=0.18U  W=1.7U  
M7      u8_G    EN      VSS     VSS     N   L=0.18U  W=0.5U  
M8      u8_G    EN      VDD     VDD     P   L=0.18U  W=1.29U  
M9      u8_S    U23_in  VSS     VSS     N   L=0.18U  W=0.42U  
M10     u8_S    U23_in  VDD     VDD     P   L=0.18U  W=1.08U  
M11     U23_in  D       VSS     VSS     N   L=0.18U  W=0.42U  
M12     U23_in  D       VDD     VDD     P   L=0.18U  W=1.08U  
M13     U26_out U26_in  VSS     VSS     N   L=0.18U  W=0.69U  
M14     U26_out U26_in  VDD     VDD     P   L=0.18U  W=1.77U  
M15     U26_in  u8_D    VSS     VSS     N   L=0.18U  W=0.69U  
M16     U26_in  u8_D    VDD     VDD     P   L=0.185U  W=1.77U  
M17     QN      u8_D    VSS     VSS     N   L=0.18U  W=2.91U  
M18     QN      u8_D    VDD     VDD     P   L=0.183U  W=8.31U  

.ENDS lanln4

.SUBCKT lanlq4 Q  D EN VDD VSS
M1      u9_S    u9_GB   u9_D    VDD     P   L=0.18U  W=1.04U    
M2      u9_S    u9_G    u9_D    VSS     N   L=0.18U  W=0.69U    
M3      U23_out u9_G    u9_S    VDD     P   L=0.18U  W=1.77U   
M4      U23_out u9_GB   u9_S    VSS     N   L=0.18U  W=0.42U    
M5      u9_G    u9_GB   VSS     VSS     N   L=0.18U  W=0.69U    
M6      u9_G    u9_GB   VDD     VDD     P   L=0.18U  W=1.73U    
M7      u9_GB   EN      VSS     VSS     N   L=0.18U  W=0.6U    
M8      u9_GB   EN      VDD     VDD     P   L=0.185U  W=1.43U    
M9      U23_out D       VSS     VSS     N   L=0.18U  W=0.42U    
M10     U23_out D       VDD     VDD     P   L=0.18U  W=1.08U    
M11     u9_D    U27_in  VSS     VSS     N   L=0.18U  W=0.69U    
M12     u9_D    U27_in  VDD     VDD     P   L=0.184U  W=1.77U    
M13     U27_in  u9_S    VSS     VSS     N   L=0.18U  W=0.69U    
M14     U27_in  u9_S    VDD     VDD     P   L=0.184U  W=1.77U    
M15     Q       u9_S    VSS     VSS     N   L=0.18U  W=2.91U    
M16     Q       u9_S    VDD     VDD     P   L=0.184U  W=8.31U    

.ENDS lanlq4

.SUBCKT mffnrb4 Q QN  CP D ENN VDD VSS
M1      u8_S    u8_GB   u8_D    VDD     P   L=0.186U  W=1.22U  
M2      u8_S    u8_G    u8_D    VSS     N   L=0.18U   W=0.47U  
M3      u9_S    u8_G    u8_S    VDD     P   L=0.18U   W=1.22U  
M4      u9_S    u8_GB   u8_S    VSS     N   L=0.18U   W=0.47U  
M5      U24_out u8_GB   U22_in  VDD     P   L=0.186U  W=1.19U  
M6      U24_out u8_G    U22_in  VSS     N   L=0.18U   W=0.47U  
M7      U27_S   U30_in  U27_D   VDD     P   L=0.18U   W=1.45U  
M8      U27_S   U30_out U27_D   VSS     N   L=0.18U   W=0.58U  
M9      U27_S   U30_out U28_D   VDD     P   L=0.18U   W=1.5U  
M10     U27_S   U30_in  U28_D   VSS     N   L=0.18U   W=0.58U  
M11     U27_S   u8_G    U22_in  VDD     P   L=0.18U   W=1.38U  
M12     U27_S   u8_GB   U22_in  VSS     N   L=0.18U   W=0.47U  
M13     u8_D    U22_in  VSS     VSS     N   L=0.18U   W=0.47U  
M14     u8_D    U22_in  VDD     VDD     P   L=0.18U   W=1.19U  
M15     U24_out u8_D    VSS     VSS     N   L=0.18U   W=0.47U  
M16     U24_out u8_D    VDD     VDD     P   L=0.18U   W=1.19U  
M17     u9_S    U23_in  VSS     VSS     N   L=0.18U   W=0.47U  
M18     u9_S    U23_in  VDD     VDD     P   L=0.186U  W=1.22U  
M19     u8_G    u8_GB   VSS     VSS     N   L=0.18U   W=0.62U  
M20     u8_G    u8_GB   VDD     VDD     P   L=0.186U  W=1.5U  
M21     u8_GB   CP      VSS     VSS     N   L=0.18U   W=0.62U  
M22     u8_GB   CP      VDD     VDD     P   L=0.18U   W=1.5U  
M23     U30_out U30_in  VSS     VSS     N   L=0.18U   W=0.58U  
M24     U30_out U30_in  VDD     VDD     P   L=0.18U   W=1.5U  
M25     U28_D   D       VSS     VSS     N   L=0.18U   W=0.58U  
M26     U28_D   D       VDD     VDD     P   L=0.186U  W=1.5U  
M27     U30_in  ENN     VSS     VSS     N   L=0.18U   W=0.58U  
M28     U30_in  ENN     VDD     VDD     P   L=0.185U  W=1.49U  
M29     U23_in  u8_S    VSS     VSS     N   L=0.18U   W=0.73U  
M30     U23_in  u8_S    VDD     VDD     P   L=0.184U  W=1.68U  
M31     Q       U23_in  VSS     VSS     N   L=0.18U   W=2.89U  
M32     Q       U23_in  VDD     VDD     P   L=0.183U  W=8.2U  
M33     QN      u8_S    VSS     VSS     N   L=0.18U   W=2.94U  
M34     QN      u8_S    VDD     VDD     P   L=0.18U   W=8.18U  
M35     U27_D   u9_S    VSS     VSS     N   L=0.18U   W=0.58U  
M36     U27_D   u9_S    VDD     VDD     P   L=0.184U  W=1.56U  

.ENDS mffnrb4

.SUBCKT mx08d1 Z  I0 I1 I2 I3 I4 I5 I6 I7 S0 S1 S2 VDD VSS
M1      i01     U102_gate U102_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M2      U47_drain U47_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M3      i01     I1      U47_drain VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M4      U103_drain S1      U102_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M5      U57_drain U47_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M6      U103_drain I3      U57_drain VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M7      U67_drain U47_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M8      U66_drain I5      U67_drain VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M9      U72_drain I7      U76_source VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M10     U76_source U47_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M11     U72_drain S1      U107_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M12     U66_drain U102_gate U107_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M13     U107_source S2      U104_source VSS     N   L=0.18U  W=0.48U   
+  PS=.300U PD=.300U
M14     U66_drain I4      U65_source VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M15     U65_source U43_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M16     U72_drain I6      U75_source VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M17     U75_source U43_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M18     i01     I0      U45_source VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M19     U45_source U43_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M20     U103_drain I2      U55_source VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M21     U55_source U43_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M22     U102_source U98_out U104_source VSS     N   L=0.18U  W=0.48U   
+  PS=.300U PD=.300U
M23     i01     I1      U42_source VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M24     U42_source U43_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M25     U53_drain U43_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M26     U103_drain I3      U53_drain VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M27     U73_drain U43_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M28     U72_drain I7      U73_drain VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M29     U66_drain I5      U62_source VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M30     U62_source U43_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M31     U61_drain U47_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M32     U66_drain I4      U61_drain VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M33     U71_drain U47_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M34     U72_drain I6      U71_drain VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M35     U41_drain U47_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M36     i01     I0      U41_drain VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M37     U51_drain U47_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M38     U103_drain I2      U51_drain VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M39     VDD     U108_gate U104_source VDD     P   L=0.18U  W=0.3U   
+  PS=.210U
M40     U43_gate S0      VSS     VSS     N   L=0.18U  W=0.69U  
M41     U43_gate S0      VDD     VDD     P   L=0.185U  W=1.45U  
M42     U102_gate S1      VSS     VSS     N   L=0.18U  W=0.42U  
M43     U102_gate S1      VDD     VDD     P   L=0.18U  W=1.11U  
M44     U98_out S2      VSS     VSS     N   L=0.18U  W=0.42U  
M45     U98_out S2      VDD     VDD     P   L=0.187U  W=1.1U  
M46     U47_gate U43_gate VSS     VSS     N   L=0.18U  W=0.51U  
M47     U47_gate U43_gate VDD     VDD     P   L=0.18U  W=1.52U  
M48     U108_gate U104_source VSS     VSS     N   L=0.18U  W=0.48U  
M49     U108_gate U104_source VDD     VDD     P   L=0.18U  W=0.24U  
M50     Z       U104_source VSS     VSS     N   L=0.18U  W=0.75U  
M51     Z       U104_source VDD     VDD     P   L=0.18U  W=1.8U  

.ENDS mx08d1

.SUBCKT mx08d2 Z  I0 I1 I2 I3 I4 I5 I6 I7 S0 S1 S2 VDD VSS
M1      U63_drain U63_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M2      U62_drain I5      U63_drain VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M3      U107_drain I7      U72_source VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M4      U72_source U63_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M5      U52_drain I3      U52_source VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M6      U52_source U63_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M7      i01     I1      U42_source VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M8      U42_source U63_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M9      U62_drain I4      U64_source VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M10     U64_source U77_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M11     U107_drain I6      U74_source VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M12     U74_source U77_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M13     U52_drain I2      U54_source VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M14     U54_source U77_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M15     U41_drain U77_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M16     i01     I0      U41_drain VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M17     VDD     U110_out U104_source VDD     P   L=0.18U  W=0.3U   
+  PS=.210U
M18     U62_drain U106_gate U106_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M19     U107_drain S1      U106_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M20     U77_drain U77_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M21     U107_drain I7      U77_drain VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M22     U62_drain I5      U66_source VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M23     U66_source U77_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M24     U52_drain I3      U56_source VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M25     U56_source U77_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M26     i01     U106_gate U102_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M27     U47_drain U77_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M28     i01     I1      U47_drain VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M29     U52_drain S1      U102_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M30     U106_source S2      U104_source VSS     N   L=0.18U  W=0.48U   
+  PS=.300U PD=.300U
M31     U78_drain U63_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M32     U107_drain I6      U78_drain VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M33     U68_drain U63_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M34     U62_drain I4      U68_drain VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M35     U58_drain U63_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M36     U52_drain I2      U58_drain VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M37     U48_drain U63_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M38     i01     I0      U48_drain VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M39     U102_source U98_out U104_source VSS     N   L=0.18U  W=0.48U   
+  PS=.300U PD=.300U
M40     U77_gate U63_gate VSS     VSS     N   L=0.18U  W=0.51U  
M41     U77_gate U63_gate VDD     VDD     P   L=0.18U  W=1.52U  
M42     U98_out S2      VSS     VSS     N   L=0.18U  W=0.42U  
M43     U98_out S2      VDD     VDD     P   L=0.187U  W=1.1U  
M44     U106_gate S1      VSS     VSS     N   L=0.18U  W=0.42U  
M45     U106_gate S1      VDD     VDD     P   L=0.18U  W=1.11U  
M46     U63_gate S0      VSS     VSS     N   L=0.18U  W=0.69U  
M47     U63_gate S0      VDD     VDD     P   L=0.185U  W=1.45U  
M48     Z       U104_source VSS     VSS     N   L=0.18U  W=1.45U  
M49     Z       U104_source VDD     VDD     P   L=0.182U  W=3.6U  
M50     U110_out U104_source VSS     VSS     N   L=0.18U  W=0.48U  
M51     U110_out U104_source VDD     VDD     P   L=0.18U  W=0.24U  

.ENDS mx08d2

.SUBCKT mx08d4 Z  I0 I1 I2 I3 I4 I5 I6 I7 S0 S1 S2 VDD VSS
M1      U63_drain U63_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M2      U62_drain I5      U63_drain VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M3      U107_drain I7      U72_source VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M4      U72_source U63_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M5      U52_drain I3      U52_source VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M6      U52_source U63_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M7      i01     I1      U42_source VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M8      U42_source U63_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M9      U62_drain I4      U64_source VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M10     U64_source U77_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M11     U107_drain I6      U74_source VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M12     U74_source U77_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M13     U52_drain I2      U54_source VDD     P   L=0.18U  W=1.47U   
+  PS=.800U PD=.800U
M14     U54_source U77_gate VDD     VDD     P   L=0.18U  W=1.47U   
+  PD=.800U
M15     U41_drain U77_gate VDD     VDD     P   L=0.18U  W=1.14U   
+  PD=.800U
M16     i01     I0      U41_drain VDD     P   L=0.18U  W=1.14U   
+  PS=.800U PD=.800U
M17     VDD     U110_out U104_source VDD     P   L=0.18U  W=0.3U   
+  PS=.210U
M18     U62_drain U106_gate U106_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M19     U107_drain S1      U106_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M20     U77_drain U77_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M21     U107_drain I7      U77_drain VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M22     U62_drain I5      U66_source VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M23     U66_source U77_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M24     U52_drain I3      U56_source VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M25     U56_source U77_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M26     i01     U106_gate U102_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M27     U47_drain U77_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M28     i01     I1      U47_drain VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M29     U52_drain S1      U102_source VSS     N   L=0.18U  W=0.47U   
+  PS=.300U PD=.433U
M30     U106_source S2      U104_source VSS     N   L=0.18U  W=0.48U   
+  PS=.300U PD=.300U
M31     U78_drain U63_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M32     U107_drain I6      U78_drain VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M33     U68_drain U63_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M34     U62_drain I4      U68_drain VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M35     U58_drain U63_gate VSS     VSS     N   L=0.18U  W=0.5U   
+  PD=.500U
M36     U52_drain I2      U58_drain VSS     N   L=0.18U  W=0.5U   
+  PS=.500U PD=.433U
M37     U48_drain U63_gate VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.500U
M38     i01     I0      U48_drain VSS     N   L=0.18U  W=0.42U   
+  PS=.500U PD=.433U
M39     U102_source U98_out U104_source VSS     N   L=0.18U  W=0.48U   
+  PS=.300U PD=.300U
M40     U77_gate U63_gate VSS     VSS     N   L=0.18U  W=0.51U  
M41     U77_gate U63_gate VDD     VDD     P   L=0.18U  W=1.52U  
M42     U98_out S2      VSS     VSS     N   L=0.18U  W=0.42U  
M43     U98_out S2      VDD     VDD     P   L=0.187U  W=1.1U  
M44     U106_gate S1      VSS     VSS     N   L=0.18U  W=0.42U  
M45     U106_gate S1      VDD     VDD     P   L=0.18U  W=1.11U  
M46     U63_gate S0      VSS     VSS     N   L=0.18U  W=0.69U  
M47     U63_gate S0      VDD     VDD     P   L=0.185U  W=1.45U  
M48     Z       U104_source VSS     VSS     N   L=0.182U  W=3U  
M49     Z       U104_source VDD     VDD     P   L=0.183U  W=7.11U  
M50     U110_out U104_source VSS     VSS     N   L=0.18U  W=0.48U  
M51     U110_out U104_source VDD     VDD     P   L=0.18U  W=0.24U  

.ENDS mx08d4

.SUBCKT nd02d7 ZN  A1 A2 VDD VSS
M1      U2_drain A2      VDD     VDD     P   L=0.18U  W=1.64U   
+  PD=1.360U
M2      U2_drain A1      VDD     VDD     P   L=0.185U  W=1.64U   
+  PD=1.360U
M3      U2_drain A1      U3_source VSS     N   L=0.18U  W=0.87U   
+  PS=.900U PD=.900U
M4      U3_source A2      VSS     VSS     N   L=0.18U  W=0.87U   
+  PD=.900U
M5      U60_out U2_drain VSS     VSS     N   L=0.18U  W=0.8U  
M6      U60_out U2_drain VDD     VDD     P   L=0.183U  W=2.26U  
M7      ZN      U60_out VSS     VSS     N   L=0.18U  W=5.12U  
M8      ZN      U60_out VDD     VDD     P   L=0.183U  W=14.34U  

.ENDS nd02d7

.SUBCKT nd02da ZN  A1 A2 VDD VSS
M1      U2_drain A2      VDD     VDD     P   L=0.18U  W=1.64U   
+  PD=1.360U
M2      U2_drain A1      VDD     VDD     P   L=0.186U  W=1.64U   
+  PD=1.360U
M3      U2_drain A1      U3_source VSS     N   L=0.18U  W=0.87U   
+  PS=.900U PD=.900U
M4      U3_source A2      VSS     VSS     N   L=0.18U  W=0.87U   
+  PD=.900U
M5      U60_out U2_drain VSS     VSS     N   L=0.18U  W=0.8U  
M6      U60_out U2_drain VDD     VDD     P   L=0.18U  W=2.26U  
M7      ZN      U60_out VSS     VSS     N   L=0.18U  W=7.14U  
M8      ZN      U60_out VDD     VDD     P   L=0.18325U  W=20.33U  

.ENDS nd02da

.SUBCKT nd03d7 ZN  A1 A2 A3 VDD VSS
M1      U5_drain A3      VDD     VDD     P   L=0.185U  W=1.29U  
M2      U5_drain A2      VDD     VDD     P   L=0.185U  W=1.29U  
M3      U5_drain A1      VDD     VDD     P   L=0.185U  W=1.29U  
M4      u2_drain A2      u2_source VSS     N   L=0.18U  W=0.83U  
M5      u2_source A3      VSS     VSS     N   L=0.18U  W=0.83U  
M6      U5_drain A1      u2_drain VSS     N   L=0.18U  W=0.83U  
M7      ZN      U34_in  VSS     VSS     N   L=0.18U  W=5.07U  
M8      ZN      U34_in  VDD     VDD     P   L=0.183U  W=14.34U  
M9      U34_in  U5_drain VSS     VSS     N   L=0.18U  W=0.8U  
M10     U34_in  U5_drain VDD     VDD     P   L=0.18U  W=2.26U  

.ENDS nd03d7

.SUBCKT nd03da ZN  A1 A2 A3 VDD VSS
M1      U5_drain A3      VDD     VDD     P   L=0.18U  W=1.29U  
M2      U5_drain A2      VDD     VDD     P   L=0.185U  W=1.29U  
M3      U5_drain A1      VDD     VDD     P   L=0.185U  W=1.29U  
M4      u2_drain A2      u2_source VSS     N   L=0.18U  W=0.83U  
M5      u2_source A3      VSS     VSS     N   L=0.18U  W=0.83U  
M6      U5_drain A1      u2_drain VSS     N   L=0.18U  W=0.83U  
M7      ZN      U34_in  VSS     VSS     N   L=0.18U  W=7.2U  
M8      ZN      U34_in  VDD     VDD     P   L=0.183125U  W=20.25U  
M9      U34_in  U5_drain VSS     VSS     N   L=0.18U  W=0.8U  
M10     U34_in  U5_drain VDD     VDD     P   L=0.18U  W=2.26U  

.ENDS nd03da

.SUBCKT nd04d7 ZN  A1 A2 A3 A4 VDD VSS
M1      U7_drain A4      VDD     VDD     P     L=0.18U   W=1.08U  
M2      U7_drain A3      VDD     VDD     P     L=0.18U   W=1.08U  
M3      U7_drain A1      VDD     VDD     P     L=0.18U   W=1.08U  
M4      U7_drain A2      VDD     VDD     P     L=0.18U   W=1.08U  
M5      U6_drain A1      U6_source VSS     N   L=0.18U   W=0.89U  
M6      U6_source A4      VSS     VSS     N    L=0.18U   W=0.89U  
M7      U7_drain A2      U4_source VSS     N   L=0.18U   W=0.89U  
M8      U4_source A3      U6_drain VSS     N   L=0.18U   W=0.89U  
M9      U33_out U7_drain VSS     VSS     N     L=0.18U   W=0.8U  
M10     U33_out U7_drain VDD     VDD     P     L=0.18U   W=2.26U  
M11     ZN      U33_out VSS     VSS     N      L=0.18U   W=5.05U  
M12     ZN      U33_out VDD     VDD     P      L=0.183U  W=14.44U  

.ENDS nd04d7

.SUBCKT nd04da ZN  A1 A2 A3 A4 VDD VSS
M1      U7_drain A4      VDD     VDD     P     L=0.18U   W=1.08U  
M2      U7_drain A3      VDD     VDD     P     L=0.18U   W=1.08U  
M3      U7_drain A1      VDD     VDD     P     L=0.18U   W=1.08U  
M4      U7_drain A2      VDD     VDD     P     L=0.18U   W=1.08U  
M5      U6_drain A1      U6_source VSS     N   L=0.18U   W=0.89U  
M6      U6_source A4      VSS     VSS     N    L=0.18U   W=0.89U  
M7      U7_drain A2      U4_source VSS     N   L=0.18U   W=0.89U  
M8      U4_source A3      U6_drain VSS     N   L=0.18U   W=0.89U  
M9      U33_out U7_drain VSS     VSS     N     L=0.18U   W=0.8U  
M10     U33_out U7_drain VDD     VDD     P     L=0.18U   W=2.26U  
M11     ZN      U33_out VSS     VSS     N      L=0.18U   W=7.14U  
M12     ZN      U33_out VDD     VDD     P      L=0.183U  W=20.33U  

.ENDS nd04da

.SUBCKT nr02d7 ZN  A1 A2 VDD VSS
M1      U36_out U36_in  VSS     VSS     N   L=0.18U  W=0.97U  
M2      U36_out U36_in  VDD     VDD     P   L=0.183U  W=2.26U  
M3      ZN      U36_out VSS     VSS     N   L=0.1865U  W=5.05U  
M4      ZN      U36_out VDD     VDD     P   L=0.18U  W=14.34U  
M5      U36_in  A1      VSS     VSS     N   L=0.18U  W=0.42U  
M6      U36_in  A2      VSS     VSS     N   L=0.18U  W=0.42U  
M7      U36_in  A2      u1_source VDD     P   L=0.187U  W=2.12U  
M8      VDD     A1      u1_source VDD     P   L=0.183U  W=2.12U  

.ENDS nr02d7

.SUBCKT nr02da ZN  A1 A2 VDD VSS
M1      U36_out U36_in  VSS     VSS     N   L=0.18U  W=0.97U  
M2      U36_out U36_in  VDD     VDD     P   L=0.183U  W=2.26U  
M3      ZN      U36_out VSS     VSS     N   L=0.18U  W=7.26U  
M4      ZN      U36_out VDD     VDD     P   L=0.182667U  W=20.3U  
M5      U36_in  A1      VSS     VSS     N   L=0.18U  W=0.42U  
M6      U36_in  A2      VSS     VSS     N   L=0.18U  W=0.42U  
M7      U36_in  A2      u1_source VDD     P   L=0.187U  W=2.12U  
M8      VDD     A1      u1_source VDD     P   L=0.183U  W=2.12U  

.ENDS nr02da

.SUBCKT nr03d7 ZN  A1 A2 A3 VDD VSS
M1      U38_drain A3      VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=1.115U
M2      U38_drain A2      VSS     VSS     N   L=0.18U  W=0.42U    
+  PD=1.115U
M3      U38_drain A1      VSS     VSS     N   L=0.18U  W=0.42U     
+  PD=1.115U
M4      U62_out U38_drain VSS     VSS     N   L=0.18U  W=0.91U    
M5      U62_out U38_drain VDD     VDD     P   L=0.184U  W=2.12U    
M6      ZN      U62_out VSS     VSS     N   L=0.183U  W=5.05U    
M7      ZN      U62_out VDD     VDD     P   L=0.182U  W=14.34U    
M8      U36_drain A3      VDD     VDD     P   L=0.184U  W=2.12U     
+  PD=1.633U
M9      U38_drain A1      u1_source VDD     P   L=0.189U  W=2.12U   
+  PS=1.595U PD=1.595U
M10     u1_source A2      U36_drain VDD     P   L=0.184U  W=2.12U     
+  PS=1.633U PD=1.595U

.ENDS nr03d7

.SUBCKT nr03da ZN  A1 A2 A3 VDD VSS
M1      U38_drain A3      VSS     VSS     N   L=0.18U  W=0.42U     
+  PD=1.115U
M2      U38_drain A2      VSS     VSS     N   L=0.18U  W=0.42U     
+  PD=1.115U
M3      U38_drain A1      VSS     VSS     N   L=0.18U  W=0.42U     
+  PD=1.115U
M4      U62_out U38_drain VSS     VSS     N   L=0.18U  W=0.9U    
M5      U62_out U38_drain VDD     VDD     P   L=0.184U  W=2.12U    
M6      ZN      U62_out VSS     VSS     N   L=0.18U  W=7.2U   
M7      ZN      U62_out VDD     VDD     P   L=0.182U  W=20.28U    
M8      U36_drain A3      VDD     VDD     P   L=0.184U  W=2.12U     
+  PD=1.633U
M9      U38_drain A1      u1_source VDD     P   L=0.188U  W=2.12U    
+  PS=1.595U PD=1.595U
M10     u1_source A2      U36_drain VDD     P   L=0.184U  W=2.12U     
+  PS=1.633U PD=1.595U

.ENDS nr03da

.SUBCKT nr04d7 ZN  A1 A2 A3 A4 VDD VSS
M1      U40_drain A4      VSS     VSS     N   L=0.18U  W=0.42U  
M2      U40_drain A3      VSS     VSS     N   L=0.18U  W=0.42U  
M3      U40_drain A2      VSS     VSS     N   L=0.18U  W=0.42U  
M4      U40_drain A1      VSS     VSS     N   L=0.18U  W=0.42U  
M5      U40_drain A1      u1_source VDD     P   L=0.185U  W=2.09U  
M6      U42_drain A3      U42_source VDD     P   L=0.18U  W=2.12U  
M7      u1_source A2      U42_drain VDD     P   L=0.18U  W=2.12U  
M8      U42_source A4      VDD     VDD     P   L=0.18U  W=2.12U  
M9      ZN      U43_in  VSS     VSS     N   L=0.184U  W=5.05U  
M10     ZN      U43_in  VDD     VDD     P   L=0.183U  W=14.34U  
M11     U43_in  U40_drain VSS     VSS     N   L=0.18U  W=1.01U  
M12     U43_in  U40_drain VDD     VDD     P   L=0.18U  W=2.26U  

.ENDS nr04d7

.SUBCKT nr04da ZN  A1 A2 A3 A4 VDD VSS
M1      U40_drain A4      VSS     VSS     N   L=0.18U  W=0.42U   
M2      U40_drain A3      VSS     VSS     N   L=0.18U  W=0.42U
M3      U40_drain A2      VSS     VSS     N   L=0.18U  W=0.42U
M4      U40_drain A1      VSS     VSS     N   L=0.18U  W=0.42U
M5      U40_drain A1      u1_source VDD     P   L=0.187U  W=2.12U
M6      U42_drain A3      U42_source VDD     P   L=0.186U  W=2.12U
M7      u1_source A2      U42_drain VDD     P   L=0.187U  W=2.12U
M8      U42_source A4      VDD     VDD     P   L=0.186U  W=2.12U
M9      ZN      U43_in  VSS     VSS     N   L=0.183U  W=7.26U
M10     ZN      U43_in  VDD     VDD     P   L=0.183U  W=20.24U
M11     U43_in  U40_drain VSS     VSS     N   L=0.18U  W=0.91U
M12     U43_in  U40_drain VDD     VDD     P   L=0.18U  W=2.4U
.ENDS nr04da

.SUBCKT or02d7 Z  A1 A2 VDD VSS
M1      u2_drain A2      VSS     VSS     N   L=0.18U    W=0.45U
+  PD=.430U
M2      Z       u2_drain VSS     VSS     N   L=0.188U   W=5.07U
+  PD=1.105U
M3      u2_drain A1      VSS     VSS     N   L=0.18U    W=0.45U
+  PD=.430U
M4      Z       u2_drain VDD     VDD     P   L=0.182U   W=14.34U
+  PD=1.380U
M5      u2_drain A1      u1_source VDD     P   L=0.187U  W=2.12U
+  PS=.840U PD=.840U
M6      VDD     A2      u1_source VDD     P   L=0.187U   W=2.12U
+  PS=.840U

.ENDS or02d7

.SUBCKT or02da Z  A1 A2 VDD VSS
M1      u2_drain A2      VSS     VSS     N   L=0.18U      W=0.45U
+  PD=.430U
M2      Z       u2_drain VSS     VSS     N   L=0.187U       W=7.2U
+  PD=1.105U
M3      u2_drain A1      VSS     VSS     N   L=0.18U      W=0.45U
+  PD=.430U
M4      Z       u2_drain VDD     VDD     P   L=0.182U      W=20.06U
+  PD=1.380U
M5      u2_drain A1      u1_source VDD     P   L=0.185U    W=2.11U
+  PS=.840U PD=.840U
M6      VDD     A2      u1_source VDD     P   L=0.186U     W=2.11U
+  PS=.840U

.ENDS or02da

.SUBCKT or03d7 Z  A1 A2 A3 VDD VSS
M1      U39_drain A3      VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.480U
M2      U39_drain A2      VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.480U
M3      U39_drain A1      VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.480U
M4      Z       U39_drain VSS     VSS     N   L=0.18U  W=5.05U  
M5      Z       U39_drain VDD     VDD     P   L=0.182U  W=14.3U  
M6      U39_drain A1      U9_source VDD     P   L=0.187U  W=2.127U   
+  PS=1.195U PD=1.195U
M7      U9_source A2      U35_source VDD     P   L=0.18U  W=2.26U   
+  PS=1.247U PD=1.195U
M8      U35_source A3      VDD     VDD     P   L=0.18U  W=2.26U   
+  PD=1.247U

.ENDS or03d7

.SUBCKT or03da Z  A1 A2 A3 VDD VSS
M1      U39_drain A3      VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.480U
M2      U39_drain A2      VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.480U
M3      U39_drain A1      VSS     VSS     N   L=0.18U  W=0.42U   
+  PD=.480U
M4      Z       U39_drain VSS     VSS     N   L=0.18U  W=7.2U  
M5      Z       U39_drain VDD     VDD     P   L=0.182U  W=20.28U  
M6      U39_drain A1      U9_source VDD     P   L=0.187U  W=2.127U   
+  PS=1.195U PD=1.195U
M7      U9_source A2      U35_source VDD     P   L=0.18U  W=2.26U   
+  PS=1.247U PD=1.195U
M8      U35_source A3      VDD     VDD     P   L=0.18U  W=2.26U   
+  PD=1.247U

.ENDS or03da

.SUBCKT or04d7 Z  A1 A2 A3 A4 VDD VSS
M1      u2_drain A2      VSS     VSS     N   L=0.18U  W=0.42U
+  PD=.450U
M2      u2_drain A3      VSS     VSS     N   L=0.18U  W=0.42U
+  PD=.450U
M3      u2_drain A4      VSS     VSS     N   L=0.18U  W=0.42U
+  PD=.450U
M4      u2_drain A1      VSS     VSS     N   L=0.18U  W=0.42U
+  PD=.450U
M5      Z       u2_drain VSS     VSS     N   L=0.18U  W=4.98U
M6      Z       u2_drain VDD     VDD     P   L=0.183U  W=14.41U
M7      U41_drain A4      VDD     VDD     P   L=0.18U  W=2.26U
+  PD=1.424U
M8      u2_drain A1      U9_source VDD     P   L=0.184U  W=2.26U
+  PS=1.410U PD=1.410U
M9      U36_drain A3      U41_drain VDD     P   L=0.18U  W=2.26U
+  PS=1.424U PD=1.410U
M10     U9_source A2      U36_drain VDD     P   L=0.183U  W=2.26U
+  PS=1.410U PD=1.410U

.ENDS or04d7

.SUBCKT or04da Z  A1 A2 A3 A4 VDD VSS
M1      u2_drain A2      VSS     VSS     N   L=0.18U  W=0.42U
+  PD=.450U
M2      u2_drain A3      VSS     VSS     N   L=0.18U  W=0.42U
+  PD=.450U
M3      u2_drain A4      VSS     VSS     N   L=0.18U  W=0.42U
+  PD=.450U
M4      u2_drain A1      VSS     VSS     N   L=0.18U  W=0.42U
+  PD=.450U
M5      Z       u2_drain VSS     VSS     N   L=0.182U  W=7.2U
M6      Z       u2_drain VDD     VDD     P   L=0.183U  W=20.28U
M7      U41_drain A4      VDD     VDD     P   L=0.18U  W=2.26U
+  PD=1.424U
M8      u2_drain A1      U9_source VDD     P   L=0.184U  W=2.26U
+  PS=1.410U PD=1.410U
M9      U36_drain A3      U41_drain VDD     P   L=0.18U  W=2.26U
+  PS=1.424U PD=1.410U
M10     U9_source A2      U36_drain VDD     P   L=0.183U  W=2.26U
+  PS=1.410U PD=1.410U

.ENDS or04da

.SUBCKT sdbfb1 Q QN  CDN CPN D SC SD SDN VDD VSS
M1      U76_out CDN     VDD     VDD     P   L=0.18U  W=1.36U  
M2      U76_out U76_in1 VDD     VDD     P   L=0.18U  W=1.36U  
M3      U76_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.79U  
M4      U76_out U76_in1 U76_$$7 VSS     N   L=0.18U  W=0.79U  
M5      U76_in1 SDN     VDD     VDD     P   L=0.18U  W=1.38U  
M6      U76_in1 U73_in1 VDD     VDD     P   L=0.186U  W=1.25U  
M7      U73_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.79U  
M8      U76_in1 U73_in1 U73_$$7 VSS     N   L=0.18U  W=0.79U  
M9      u9_S    SDN     VDD     VDD     P   L=0.186U  W=1.38U  
M10     u9_S    U74_in1 VDD     VDD     P   L=0.18U  W=1.38U  
M11     U74_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.83U  
M12     u9_S    U74_in1 U74_$$7 VSS     N   L=0.18U  W=0.83U  
M13     U74_in1 CDN     VDD     VDD     P   L=0.186U  W=1.38U  
M14     U74_in1 u9_D    VDD     VDD     P   L=0.186U  W=1.38U  
M15     U75_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.83U  
M16     U74_in1 u9_D    U75_$$7 VSS     N   L=0.18U  W=0.83U  
M17     U66_drain SD      U66_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M18     VDD     U45_gate U66_drain VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M19     U67_drain D       U66_source VDD     P   L=0.185U  W=1.78U   
+  PS=.520U PD=.520U
M20     VDD     U43_gate U67_drain VDD     P   L=0.185U  W=1.78U   
+  PS=.520U
M21     U68_drain U45_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M22     U66_source D       U68_drain VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M23     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U   
+  PD=.480U
M24     U66_source SD      U69_drain VSS     N   L=0.18U  W=0.66U   
+  PS=.480U PD=.480U
M25     U76_out u7_GB   U73_in1 VDD     P   L=0.187U  W=1.25U  
M26     U76_out u7_G    U73_in1 VSS     N   L=0.18U  W=0.46U  
M27     U66_source u7_G    U73_in1 VDD     P   L=0.186U  W=1.25U   
+  PD=.520U
M28     U66_source u7_GB   U73_in1 VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M29     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.73U  
M30     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M31     U76_in1 u7_GB   u9_D    VDD     P   L=0.18U  W=0.73U  
M32     U76_in1 u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  
M33     u7_G    CPN     VSS     VSS     N   L=0.18U  W=0.69U  
M34     u7_G    CPN     VDD     VDD     P   L=0.184U  W=1.8U  
M35     u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.69U  
M36     u7_GB   u7_G    VDD     VDD     P   L=0.184U  W=1.8U  
M37     U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M38     U43_gate U45_gate VDD     VDD     P   L=0.184U  W=1.91U  
M39     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M40     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M41     QN      u9_D    VSS     VSS     N   L=0.18U  W=0.69U  
M42     QN      u9_D    VDD     VDD     P   L=0.184U  W=1.86U  
M43     Q       U74_in1 VSS     VSS     N   L=0.18U  W=0.69U  
M44     Q       U74_in1 VDD     VDD     P   L=0.184U  W=1.86U  

.ENDS sdbfb1

.SUBCKT sdbfb2 Q QN  CDN CPN D SC SD SDN VDD VSS
M1      U76_out CDN     VDD     VDD     P   L=0.18U      W=1.36U
M2      U76_out U76_in1 VDD     VDD     P   L=0.18U      W=1.36U
M3      U76_$$7 CDN     VSS     VSS     N   L=0.18U      W=0.79U
M4      U76_out U76_in1 U76_$$7 VSS     N   L=0.18U      W=0.79U
M5      U76_in1 SDN     VDD     VDD     P   L=0.18U      W=1.38U
M6      U76_in1 U73_in1 VDD     VDD     P   L=0.186U      W=1.25U
M7      U73_$$7 SDN     VSS     VSS     N   L=0.18U      W=0.79U
M8      U76_in1 U73_in1 U73_$$7 VSS     N   L=0.18U      W=0.79U
M9      u9_S    SDN     VDD     VDD     P   L=0.186U      W=1.38U
M10     u9_S    U74_in1 VDD     VDD     P   L=0.18U      W=1.38U
M11     U74_$$7 SDN     VSS     VSS     N   L=0.18U      W=0.83U
M12     u9_S    U74_in1 U74_$$7 VSS     N   L=0.18U      W=0.83U
M13     U74_in1 CDN     VDD     VDD     P   L=0.186U      W=1.38U
M14     U74_in1 u9_D    VDD     VDD     P   L=0.186U      W=1.38U
M15     U75_$$7 CDN     VSS     VSS     N   L=0.18U      W=0.83U
M16     U74_in1 u9_D    U75_$$7 VSS     N   L=0.18U      W=0.83U
M17     U66_drain SD      U66_source VDD     P   L=0.18U       W=1.91U
+  PS=.520U PD=.520U
M18     VDD     U45_gate U66_drain VDD     P   L=0.18U       W=1.91U
+  PS=.520U
M19     U67_drain D       U66_source VDD     P   L=0.185U       W=1.78U
+  PS=.520U PD=.520U
M20     VDD     U43_gate U67_drain VDD     P   L=0.185U       W=1.78U
+  PS=.520U
M21     U68_drain U45_gate VSS     VSS     N   L=0.18U       W=0.69U
+  PD=.480U
M22     U66_source D       U68_drain VSS     N   L=0.18U       W=0.69U
+  PS=.480U PD=.480U
M23     U69_drain U43_gate VSS     VSS     N   L=0.18U       W=0.66U
+  PD=.480U
M24     U66_source SD      U69_drain VSS     N   L=0.18U       W=0.66U
+  PS=.480U PD=.480U
M25     U76_out u7_GB   U73_in1 VDD     P   L=0.185U      W=1.25U
M26     U76_out u7_G    U73_in1 VSS     N   L=0.18U      W=0.46U
M27     U66_source u7_G    U73_in1 VDD     P   L=0.18U       W=1.25U
+  PD=.520U
M28     U66_source u7_GB   U73_in1 VSS     N   L=0.18U       W=0.46U
+  PD=.480U
M29     u9_S    u7_G    u9_D    VDD     P   L=0.18U      W=0.73U
M30     u9_S    u7_GB   u9_D    VSS     N   L=0.18U      W=0.42U
M31     U76_in1 u7_GB   u9_D    VDD     P   L=0.18U      W=0.73U
M32     U76_in1 u7_G    u9_D    VSS     N   L=0.18U      W=0.46U
M33     u7_G    CPN     VSS     VSS     N   L=0.18U      W=0.69U
M34     u7_G    CPN     VDD     VDD     P   L=0.184U      W=1.8U
M35     u7_GB   u7_G    VSS     VSS     N   L=0.18U      W=0.69U
M36     u7_GB   u7_G    VDD     VDD     P   L=0.184U      W=1.8U
M37     U43_gate U45_gate VSS     VSS     N   L=0.18U      W=0.69U
M38     U43_gate U45_gate VDD     VDD     P   L=0.18U      W=1.91U
M39     U45_gate SC      VSS     VSS     N   L=0.18U      W=0.69U
M40     U45_gate SC      VDD     VDD     P   L=0.184U      W=1.91U
M41     Q       U74_in1 VSS     VSS     N   L=0.18U      W=1.5U
M42     Q       U74_in1 VDD     VDD     P   L=0.184U      W=4.1U
M43     QN      u9_D    VSS     VSS     N   L=0.18U      W=1.5U
M44     QN      u9_D    VDD     VDD     P   L=0.184U      W=4.1U

.ENDS sdbfb2

.SUBCKT sdbfb4 Q QN  CDN CPN D SC SD SDN VDD VSS
M1      U76_out CDN     VDD     VDD     P   L=0.18U  W=1.36U  
M2      U76_out U76_in1 VDD     VDD     P   L=0.18U  W=1.36U  
M3      U76_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.79U  
M4      U76_out U76_in1 U76_$$7 VSS     N   L=0.18U  W=0.79U  
M5      U76_in1 SDN     VDD     VDD     P   L=0.18U  W=1.38U  
M6      U76_in1 U73_in1 VDD     VDD     P   L=0.186U  W=1.25U  
M7      U73_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.79U  
M8      U76_in1 U73_in1 U73_$$7 VSS     N   L=0.18U  W=0.79U  
M9      u9_S    SDN     VDD     VDD     P   L=0.186U  W=1.38U  
M10     u9_S    U74_in1 VDD     VDD     P   L=0.18U  W=1.38U  
M11     U74_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.83U  
M12     u9_S    U74_in1 U74_$$7 VSS     N   L=0.18U  W=0.83U  
M13     U74_in1 CDN     VDD     VDD     P   L=0.186U  W=1.38U  
M14     U74_in1 u9_D    VDD     VDD     P   L=0.186U  W=1.38U  
M15     U75_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.83U  
M16     U74_in1 u9_D    U75_$$7 VSS     N   L=0.18U  W=0.83U  
M17     U66_drain SD      U66_source VDD     P   L=0.18U  W=1.91U   
+  PS=.520U PD=.520U
M18     VDD     U45_gate U66_drain VDD     P   L=0.18U  W=1.91U   
+  PS=.520U
M19     U67_drain D       U66_source VDD     P   L=0.185U  W=1.78U   
+  PS=.520U PD=.520U
M20     VDD     U43_gate U67_drain VDD     P   L=0.185U  W=1.78U   
+  PS=.520U
M21     U68_drain U45_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M22     U66_source D       U68_drain VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M23     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U   
+  PD=.480U
M24     U66_source SD      U69_drain VSS     N   L=0.18U  W=0.66U   
+  PS=.480U PD=.480U
M25     U76_out u7_GB   U73_in1 VDD     P   L=0.187U  W=1.25U  
M26     U76_out u7_G    U73_in1 VSS     N   L=0.18U  W=0.46U  
M27     U66_source u7_G    U73_in1 VDD     P   L=0.18U  W=1.25U   
+  PD=.520U
M28     U66_source u7_GB   U73_in1 VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M29     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.73U  
M30     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M31     U76_in1 u7_GB   u9_D    VDD     P   L=0.18U  W=0.73U  
M32     U76_in1 u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  
M33     u7_G    CPN     VSS     VSS     N   L=0.18U  W=0.69U  
M34     u7_G    CPN     VDD     VDD     P   L=0.184U  W=1.8U  
M35     u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.69U  
M36     u7_GB   u7_G    VDD     VDD     P   L=0.184U  W=1.8U  
M37     U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M38     U43_gate U45_gate VDD     VDD     P   L=0.18U  W=1.91U  
M39     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M40     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M41     Q       U74_in1 VSS     VSS     N   L=0.18U  W=2.88U  
M42     Q       U74_in1 VDD     VDD     P   L=0.184U  W=8.2U  
M43     QN      u9_D    VSS     VSS     N   L=0.18U  W=2.88U  
M44     QN      u9_D    VDD     VDD     P   L=0.184U  W=8.2U  

.ENDS sdbfb4

.SUBCKT sdbrb4 Q QN  CDN CP D SC SD SDN VDD VSS
M1      U76_out CDN     VDD     VDD     P   L=0.18U  W=1.36U  
M2      U76_out U76_in1 VDD     VDD     P   L=0.18U  W=1.36U  
M3      U76_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.79U  
M4      U76_out U76_in1 U76_$$7 VSS     N   L=0.18U  W=0.79U  
M5      U76_in1 SDN     VDD     VDD     P   L=0.18U  W=1.38U  
M6      U76_in1 U73_in1 VDD     VDD     P   L=0.186U  W=1.25U  
M7      U73_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.79U  
M8      U76_in1 U73_in1 U73_$$7 VSS     N   L=0.18U  W=0.79U  
M9      U74_out SDN     VDD     VDD     P   L=0.186U  W=1.38U  
M10     U74_out U74_in1 VDD     VDD     P   L=0.18U  W=1.38U  
M11     U74_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.83U
M12     U74_out U74_in1 U74_$$7 VSS     N   L=0.18U  W=0.83U  
M13     U74_in1 CDN     VDD     VDD     P   L=0.186U  W=1.38U  
M14     U74_in1 u9_D    VDD     VDD     P   L=0.186U  W=1.38U  
M15     U75_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.83U  
M16     U74_in1 u9_D    U75_$$7 VSS     N   L=0.18U  W=0.83U  
M17     U66_drain SD      U66_source VDD     P   L=0.18U  W=1.91U   
+  PS=.520U PD=.520U
M18     VDD     U45_gate U66_drain VDD     P   L=0.18U  W=1.91U   
+  PS=.520U
M19     VDD     U43_gate U43_source VDD     P   L=0.185U  W=1.78U   
+  PS=.520U
M20     U43_source D       U66_source VDD     P   L=0.185U  W=1.78U   
+  PS=.520U PD=.520U
M21     U68_drain U45_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M22     U66_source D       U68_drain VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M23     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U   
+  PD=.480U
M24     U66_source SD      U69_drain VSS     N   L=0.18U  W=0.66U   
+  PS=.480U PD=.480U
M25     U76_out u7_GB   U73_in1 VDD     P   L=0.187U  W=1.25U  
M26     U76_out u7_G    U73_in1 VSS     N   L=0.18U  W=0.46U  
M27     U66_source u7_G    U73_in1 VDD     P   L=0.18U  W=1.25U   
+  PD=.520U
M28     U66_source u7_GB   U73_in1 VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M29     U74_out u7_G    u9_D    VDD     P   L=0.18U  W=0.73U  
M30     U74_out u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M31     U76_in1 u7_GB   u9_D    VDD     P   L=0.18U  W=0.73U  
M32     U76_in1 u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  
M33     u7_GB   CP      VSS     VSS     N   L=0.18U  W=0.69U  
M34     u7_GB   CP      VDD     VDD     P   L=0.184U  W=1.8U  
M35     u7_G    u7_GB   VSS     VSS     N   L=0.18U  W=0.69U  
M36     u7_G    u7_GB   VDD     VDD     P   L=0.184U  W=1.8U  
M37     U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M38     U43_gate U45_gate VDD     VDD     P   L=0.18U  W=1.91U  
M39     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M40     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M41     Q       U74_in1 VSS     VSS     N   L=0.18U  W=2.99U  
M42     Q       U74_in1 VDD     VDD     P   L=0.184U  W=8.2U  
M43     QN      u9_D    VSS     VSS     N   L=0.18U  W=2.99U  
M44     QN      u9_D    VDD     VDD     P   L=0.184U  W=8.2U  

.ENDS sdbrb4

.SUBCKT sdcfb1 Q QN  CDN CPN D SC SD VDD VSS
M1      U77_out U77_in  VSS     VSS     N     L=0.18U     W=0.79U  
M2      U77_out U77_in  VDD     VDD     P     L=0.184U    W=1.73U  
M3      U15_GB  CPN     VSS     VSS     N     L=0.18U     W=0.69U  
M4      U15_GB  CPN     VDD     VDD     P     L=0.184U    W=1.81U  
M5      U15_G   U15_GB  VSS     VSS     N     L=0.18U     W=0.69U  
M6      U15_G   U15_GB  VDD     VDD     P     L=0.184U    W=1.81U  
M7      U43_gate U45_gate VSS     VSS     N   L=0.18U     W=0.69U  
M8      U43_gate U45_gate VDD     VDD     P   L=0.184U    W=1.91U  
M9      U45_gate SC      VSS     VSS     N    L=0.18U     W=0.69U  
M10     U45_gate SC      VDD     VDD     P    L=0.184U    W=1.91U  
M11     u9_S    U78_in  VSS     VSS     N     L=0.18U     W=0.83U  
M12     u9_S    U78_in  VDD     VDD     P     L=0.184U    W=1.84U  
M13     QN      u8_D    VSS     VSS     N     L=0.18U     W=0.69U  
M14     QN      u8_D    VDD     VDD     P     L=0.184U    W=2.05U  
M15     Q       U78_in  VSS     VSS     N     L=0.18U     W=0.69U  
M16     Q       U78_in  VDD     VDD     P     L=0.184U    W=2.05U  
M17     U76_out CDN     VDD     VDD     P     L=0.186U    W=1.36U  
M18     U76_out U77_out VDD     VDD     P     L=0.18U     W=1.36U  
M19     U76_$$7 CDN     VSS     VSS     N     L=0.18U     W=0.79U  
M20     U76_out U77_out U76_$$7 VSS     N     L=0.18U     W=0.79U  
M21     U78_in  CDN     VDD     VDD     P     L=0.186U     W=1.38U  
M22     U78_in  u8_D    VDD     VDD     P     L=0.18U     W=1.38U  
M23     U75_$$7 CDN     VSS     VSS     N     L=0.18U     W=0.83U  
M24     U78_in  u8_D    U75_$$7 VSS     N     L=0.18U     W=0.83U  
M25     U15_S   U15_GB  U77_in  VDD     P     L=0.18U     W=1.25U   PD=.520U
M26     U15_S   U15_G   U77_in  VSS     N     L=0.18U     W=0.46U   PD=.480U
M27     U76_out U15_G   U77_in  VDD     P     L=0.19U     W=1.25U  
M28     U76_out U15_GB  U77_in  VSS     N     L=0.18U     W=0.46U  
M29     U77_out U15_G   u8_D    VDD     P     L=0.18U     W=1.12U  
M30     U77_out U15_GB  u8_D    VSS     N     L=0.18U     W=0.46U  
M31     u9_S    U15_GB  u8_D    VDD     P     L=0.186U    W=1.12U  
M32     u9_S    U15_G   u8_D    VSS     N     L=0.18U     W=0.42U  
M33     VDD     U43_gate U43_source VDD   P   L=0.185U    W=1.78U   
+  PS=.520U
M34     U43_source D       U15_S   VDD    P   L=0.185U    W=1.78U   
+  PS=.520U PD=.520U
M35     U66_drain SD      U15_S   VDD     P   L=0.184U    W=1.91U   
+  PS=.520U PD=.520U
M36     VDD     U45_gate U66_drain VDD    P   L=0.184U    W=1.91U   
+  PS=.520U
M37     U68_drain U45_gate VSS     VSS    N   L=0.18U     W=0.69U   
+  PD=.480U
M38     U69_drain U43_gate VSS     VSS    N   L=0.18U     W=.66U   
+  PD=.480U
M39     U15_S   D       U68_drain VSS     N   L=0.18U     W=0.69U   
+  PS=.480U PD=.480U
M40     U15_S   SD      U69_drain VSS     N   L=0.18U     W=0.66U   
+  PS=.480U PD=.480U

.ENDS sdcfb1

.SUBCKT sdcfb2 Q QN  CDN CPN D SC SD VDD VSS
M1      U77_out U77_in  VSS     VSS       N   L=0.18U     W=0.79U  
M2      U77_out U77_in  VDD     VDD       P   L=0.184U    W=1.73U  
M3      U15_GB  CPN     VSS     VSS       N   L=0.18U     W=0.69U  
M4      U15_GB  CPN     VDD     VDD       P   L=0.184U    W=1.8U  
M5      U15_G   U15_GB  VSS     VSS       N   L=0.18U     W=0.69U  
M6      U15_G   U15_GB  VDD     VDD       P   L=0.184U    W=1.84U  
M7      U43_gate U45_gate VSS     VSS     N   L=0.18U     W=0.69U  
M8      U43_gate U45_gate VDD     VDD     P   L=0.184U    W=1.91U  
M9      U45_gate SC      VSS     VSS      N   L=0.18U     W=0.69U  
M10     U45_gate SC      VDD     VDD      P   L=0.184U    W=1.91U  
M11     u9_S    U78_in  VSS     VSS       N   L=0.18U     W=0.83U  
M12     u9_S    U78_in  VDD     VDD       P   L=0.184U    W=1.84U  
M13     QN      u8_D    VSS     VSS       N   L=0.18U     W=1.38U  
M14     QN      u8_D    VDD     VDD       P   L=0.182U    W=4.1U  
M15     Q       U78_in  VSS     VSS       N   L=0.18U     W=1.44U  
M16     Q       U78_in  VDD     VDD       P   L=0.184U    W=4.1U  
M17     U76_out CDN     VDD     VDD       P   L=0.186U    W=1.36U  
M18     U76_out U77_out VDD     VDD       P   L=0.18U     W=1.36U  
M19     U76_$$7 CDN     VSS     VSS       N   L=0.18U     W=0.79U  
M20     U76_out U77_out U76_$$7 VSS       N   L=0.18U     W=0.79U  
M21     U78_in  CDN     VDD     VDD       P   L=0.186U    W=1.38U  
M22     U78_in  u8_D    VDD     VDD       P   L=0.18U     W=1.38U  
M23     U75_$$7 CDN     VSS     VSS       N   L=0.18U     W=0.83U  
M24     U78_in  u8_D    U75_$$7 VSS       N   L=0.18U     W=0.83U  
M25     U15_S   U15_GB  U77_in  VDD       P   L=0.18U     W=1.25U   PD=.520U
M26     U15_S   U15_G   U77_in  VSS       N   L=0.18U     W=0.46U   PD=.480U
M27     U76_out U15_G   U77_in  VDD       P   L=0.19U     W=1.25U  
M28     U76_out U15_GB  U77_in  VSS       N   L=0.18U     W=0.46U  
M29     U77_out U15_G   u8_D    VDD       P   L=0.18U     W=1.12U  
M30     U77_out U15_GB  u8_D    VSS       N   L=0.18U     W=0.46U  
M31     u9_S    U15_GB  u8_D    VDD       P   L=0.186U    W=1.12U  
M32     u9_S    U15_G   u8_D    VSS       N   L=0.18U     W=0.42U  
M33     VDD     U43_gate U43_source VDD   P   L=0.185U    W=1.78U   
+  PS=.520U
M34     U43_source D       U15_S   VDD    P   L=0.185U    W=1.78U   
+  PS=.520U PD=.520U
M35     U66_drain SD      U15_S   VDD     P   L=0.184U    W=1.91U   
+  PS=.520U PD=.520U
M36     VDD     U45_gate U66_drain VDD    P   L=0.184U    W=1.91U   
+  PS=.520U
M37     U68_drain U45_gate VSS     VSS    N   L=0.18U     W=0.69U   
+  PD=.480U
M38     U69_drain U43_gate VSS     VSS    N   L=0.18U     W=.66U   
+  PD=.480U
M39     U15_S   D       U68_drain VSS     N   L=0.18U     W=0.69U   
+  PS=.480U PD=.480U
M40     U15_S   SD      U69_drain VSS     N   L=0.18U     W=.66U   
+  PS=.480U PD=.480U

.ENDS sdcfb2

.SUBCKT sdcfb4 Q QN  CDN CPN D SC SD VDD VSS
M1      U77_out U77_in  VSS     VSS     N        L=0.18U     W=0.79U  
M2      U77_out U77_in  VDD     VDD     P        L=0.184U    W=1.73U  
M3      U15_GB  CPN     VSS     VSS     N        L=0.18U     W=0.69U  
M4      U15_GB  CPN     VDD     VDD     P        L=0.186U    W=1.8U  
M5      U15_G   U15_GB  VSS     VSS     N        L=0.18U     W=0.69U  
M6      U15_G   U15_GB  VDD     VDD     P        L=0.184U    W=1.8U  
M7      U43_gate U45_gate VSS     VSS     N      L=0.18U     W=0.69U  
M8      U43_gate U45_gate VDD     VDD     P      L=0.184U    W=1.91U  
M9      U45_gate SC      VSS     VSS     N       L=0.18U     W=0.69U  
M10     U45_gate SC      VDD     VDD     P       L=0.184U    W=1.91U  
M11     u9_S    U78_in  VSS     VSS     N        L=0.18U     W=0.83U  
M12     u9_S    U78_in  VDD     VDD     P        L=0.184U    W=1.84U  
M13     QN      u8_D    VSS     VSS     N        L=0.18U     W=2.88U  
M14     QN      u8_D    VDD     VDD     P        L=0.184U    W=8.2U  
M15     Q       U78_in  VSS     VSS     N        L=0.184U    W=2.88U  
M16     Q       U78_in  VDD     VDD     P        L=0.185U    W=8.2U  
M17     U76_out CDN     VDD     VDD     P        L=0.186U    W=1.36U  
M18     U76_out U77_out VDD     VDD     P        L=0.18U     W=1.36U  
M19     U76_$$7 CDN     VSS     VSS     N        L=0.18U     W=0.69U  
M20     U76_out U77_out U76_$$7 VSS     N        L=0.18U     W=0.69U  
M21     U78_in  CDN     VDD     VDD     P        L=0.186U    W=1.38U  
M22     U78_in  u8_D    VDD     VDD     P        L=0.18U     W=1.38U  
M23     U75_$$7 CDN     VSS     VSS     N        L=0.18U     W=0.83U  
M24     U78_in  u8_D    U75_$$7 VSS     N        L=0.18U     W=0.83U  
M25     U15_S   U15_GB  U77_in  VDD     P        L=0.18U     W=1.25U   PD=.520U
M26     U15_S   U15_G   U77_in  VSS     N        L=0.18U     W=0.46U   PD=.480U
M27     U76_out U15_G   U77_in  VDD     P        L=0.186U    W=1.25U  
M28     U76_out U15_GB  U77_in  VSS     N        L=0.18U     W=0.46U  
M29     U77_out U15_G   u8_D    VDD     P        L=0.18U     W=1.12U  
M30     U77_out U15_GB  u8_D    VSS     N        L=0.18U     W=0.46U  
M31     u9_S    U15_GB  u8_D    VDD     P        L=0.186U    W=1.12U  
M32     u9_S    U15_G   u8_D    VSS     N        L=0.18U     W=0.42U  
M33     VDD     U43_gate U43_source VDD     P    L=0.185U    W=1.78U   
+  PS=.520U
M34     U43_source D       U15_S   VDD     P     L=0.185U    W=1.78U   
+  PS=.520U PD=.520U
M35     U66_drain SD      U15_S   VDD     P      L=0.184U    W=1.91U   
+  PS=.520U PD=.520U
M36     VDD     U45_gate U66_drain VDD     P     L=0.184U    W=1.91U   
+  PS=.520U
M37     U68_drain U45_gate VSS     VSS     N     L=0.18U     W=0.69U   
+  PD=.480U
M38     U69_drain U43_gate VSS     VSS     N     L=0.18U     W=.66U   
+  PD=.480U
M39     U15_S   D       U68_drain VSS     N      L=0.18U     W=0.69U   
+  PS=.480U PD=.480U
M40     U15_S   SD      U69_drain VSS     N      L=0.18U     W=.66U   
+  PS=.480U PD=.480U

.ENDS sdcfb4

.SUBCKT sdcfq4 Q  CDN CPN D SC SD VDD VSS
M1      U77_out U77_in  VSS     VSS     N   L=0.18U     W=0.82U
M2      U77_out U77_in  VDD     VDD     P   L=0.185U    W=1.66U
M3      U15_GB  CPN     VSS     VSS     N   L=0.18U    W=0.66U
M4      U15_GB  CPN     VDD     VDD     P   L=0.185U     W=1.74U
M5      U15_G   U15_GB  VSS     VSS     N   L=0.18U     W=0.66U
M6      U15_G   U15_GB  VDD     VDD     P   L=0.184U    W=1.74U
M7      U43_gate U45_gate VSS     VSS     N   L=0.18U    W=0.69U
M8      U43_gate U45_gate VDD     VDD     P   L=0.18U      W=1.91U
M9      U45_gate SC      VSS     VSS     N   L=0.18U    W=0.69U
M10     U45_gate SC      VDD     VDD     P   L=0.184U    W=1.91U
M11     U78_out U78_in  VSS     VSS     N   L=0.18U     W=0.83U
M12     U78_out U78_in  VDD     VDD     P   L=0.18U   W=1.66U
M13     Q       U78_in  VSS     VSS     N   L=0.1823333U    W=2.88U
M14     Q       U78_in  VDD     VDD     P   L=0.18225U    W=8.2U
M15     U76_out CDN     VDD     VDD     P   L=0.186U     W=1.36U
M16     U76_out U77_out VDD     VDD     P   L=0.186U     W=1.36U
M17     U76_$$7 CDN     VSS     VSS     N   L=0.18U    W=0.82U
M18     U76_out U77_out U76_$$7 VSS     N   L=0.18U    W=0.82U
M19     U78_in  CDN     VDD     VDD     P   L=0.185U      W=1.45U
M20     U78_in  u8_D    VDD     VDD     P   L=0.185U    W=1.45U
M21     U75_$$7 CDN     VSS     VSS     N   L=0.18U     W=0.83U
M22     U78_in  u8_D    U75_$$7 VSS     N   L=0.18U      W=0.83U
M23     VDD     U45_gate U45_source VDD     P   L=0.18U       W=1.91U
+  PS=.520U
M24     VDD     U43_gate U43_source VDD     P   L=0.184U      W=1.78U
+  PS=.520U
M25     U43_source D       U15_S   VDD     P   L=0.184U       W=1.78U
+  PS=.520U PD=.520U
M26     U45_source SD      U15_S   VDD     P   L=0.18U    W=1.91U
+  PS=.520U PD=.520U
M27     U15_S   U15_GB  U77_in  VDD     P   L=0.186U    PD=.520U  W=1.38U
M28     U15_S   U15_G   U77_in  VSS     N   L=0.18U    PD=.480U  W=0.42U
M29     U76_out U15_G   U77_in  VDD     P   L=0.186U      W=1.38U
M30     U76_out U15_GB  U77_in  VSS     N   L=0.18U     W=0.46U
M31     U77_out U15_G   u8_D    VDD     P   L=0.18U    W=0.69U
M32     U77_out U15_GB  u8_D    VSS     N   L=0.18U     W=0.46U
M33     U78_out U15_GB  u8_D    VDD     P   L=0.18U     W=0.69U
M34     U78_out U15_G   u8_D    VSS     N   L=0.18U    W=0.46U
M35     U68_drain U45_gate VSS     VSS     N   L=0.18U   W=0.69U
+  PD=.480U
M36     U69_drain U43_gate VSS     VSS     N   L=0.18U    W=0.66U
+  PD=.480U
M37     U15_S   SD      U69_drain VSS     N   L=0.18U   W=0.66U
+  PS=.480U PD=.480U
M38     U15_S   D       U68_drain VSS     N   L=0.18U    W=0.69U
+  PS=.480U PD=.480U

.ENDS sdcfq4

.SUBCKT sdcrb4 Q QN  CDN CP D SC SD VDD VSS
M1      U77_out U77_in  VSS     VSS     N   L=0.18U     W=0.82U
M2      U77_out U77_in  VDD     VDD     P   L=0.185U    W=1.66U
M3      U15_G   CP      VSS     VSS     N   L=0.18U     W=0.66U
M4      U15_G   CP      VDD     VDD     P   L=0.184U    W=1.74U
M5      U15_GB  U15_G   VSS     VSS     N   L=0.18U     W=0.66U
M6      U15_GB  U15_G   VDD     VDD     P   L=0.18U   W=1.74U
M7      U43_gate U45_gate VSS     VSS     N   L=0.18U    W=0.69U
M8      U43_gate U45_gate VDD     VDD     P   L=0.18U    W=1.91U
M9      U45_gate SC      VSS     VSS     N   L=0.18U   W=0.69U
M10     U45_gate SC      VDD     VDD     P   L=0.184U    W=1.91U
M11     u9_S    U78_in  VSS     VSS     N   L=0.18U    W=0.83U
M12     u9_S    U78_in  VDD     VDD     P   L=0.185U      W=1.66U
M13     QN      u8_D    VSS     VSS     N   L=0.18U     W=2.95U
M14     QN      u8_D    VDD     VDD     P   L=0.183U     W=8.2U
M15     Q       U78_in  VSS     VSS     N   L=0.18U     W=2.95U
M16     Q       U78_in  VDD     VDD     P   L=0.182U     W=8.2U
M17     U76_out CDN     VDD     VDD     P   L=0.186U    W=1.36U
M18     U76_out U77_out VDD     VDD     P   L=0.18U    W=1.36U
M19     U76_$$7 CDN     VSS     VSS     N   L=0.18U     W=0.82U
M20     U76_out U77_out U76_$$7 VSS     N   L=0.18U    W=0.82U
M21     U78_in  CDN     VDD     VDD     P   L=0.185U    W=1.45U
M22     U78_in  u8_D    VDD     VDD     P   L=0.18U    W=1.45U
M23     U75_$$7 CDN     VSS     VSS     N   L=0.18U    W=0.83U
M24     U78_in  u8_D    U75_$$7 VSS     N   L=0.18U    W=0.83U
M25     U15_S   U15_GB  U77_in  VDD     P   L=0.18U  PD=.520U  W=1.38U
M26     U15_S   U15_G   U77_in  VSS     N   L=0.18U  PD=.480U  W=0.42U
M27     U76_out U15_G   U77_in  VDD     P   L=0.186U  W=1.38U
M28     U76_out U15_GB  U77_in  VSS     N   L=0.18U    W=0.46U
M29     U77_out U15_G   u8_D    VDD     P   L=0.18U    W=0.69U
M30     U77_out U15_GB  u8_D    VSS     N   L=0.18U   W=0.46U
M31     u9_S    U15_GB  u8_D    VDD     P   L=0.18U     W=0.69U
M32     u9_S    U15_G   u8_D    VSS     N   L=0.18U    W=0.42U
M33     U67_drain D       U15_S   VDD     P   L=0.184U    W=1.78U
+  PS=.520U PD=.520U
M34     VDD     U43_gate U67_drain VDD     P   L=0.184U   W=1.78U
+  PS=.520U
M35     U66_drain SD      U15_S   VDD     P   L=0.18U     W=1.91U
+  PS=.520U PD=.520U
M36     VDD     U45_gate U66_drain VDD     P   L=0.18U     W=1.91U
+  PS=.520U
M37     U68_drain U45_gate VSS     VSS     N   L=0.18U    W=0.69U
+  PD=.480U
M38     U69_drain U43_gate VSS     VSS     N   L=0.18U   W=0.66U
+  PD=.480U
M39     U15_S   D       U68_drain VSS     N   L=0.18U   W=0.69U
+  PS=.480U PD=.480U
M40     U15_S   SD      U69_drain VSS     N   L=0.18U    W=0.66U
+  PS=.480U PD=.480U

.ENDS sdcrb4

.SUBCKT sdcrn4 QN  CDN CP D SC SD VDD VSS
M1      U77_out U77_in  VSS     VSS     N      L=0.18U     W=0.82U  
M2      U77_out U77_in  VDD     VDD     P      L=0.185U    W=1.66U  
M3      U15_G   CP      VSS     VSS     N      L=0.18U     W=0.66U  
M4      U15_G   CP      VDD     VDD     P      L=0.18U     W=1.74U  
M5      U15_GB  U15_G   VSS     VSS     N      L=0.18U     W=0.66U  
M6      U15_GB  U15_G   VDD     VDD     P      L=0.184U    W=1.74U  
M7      U43_gate U45_gate VSS     VSS     N    L=0.18U     W=0.69U  
M8      U43_gate U45_gate VDD     VDD     P    L=0.184U    W=1.91U  
M9      U45_gate SC      VSS     VSS     N     L=0.18U     W=0.69U  
M10     U45_gate SC      VDD     VDD     P     L=0.184U    W=1.91U  
M11     u9_S    U78_in  VSS     VSS     N      L=0.18U     W=0.83U  
M12     u9_S    U78_in  VDD     VDD     P      L=0.184U    W=1.66U  
M13     QN      u8_D    VSS     VSS     N      L=0.18U     W=2.88U  
M14     QN      u8_D    VDD     VDD     P      L=0.184U    W=8.2U  
M15     U76_out CDN     VDD     VDD     P      L=0.186U    W=1.36U  
M16     U76_out U77_out VDD     VDD     P      L=0.18U     W=1.36U  
M17     U76_$$7 CDN     VSS     VSS     N      L=0.18U     W=0.82U  
M18     U76_out U77_out U76_$$7 VSS     N      L=0.18U     W=0.82U  
M19     U78_in  CDN     VDD     VDD     P      L=0.185U    W=1.45U  
M20     U78_in  u8_D    VDD     VDD     P      L=0.18U     W=1.45U  
M21     U75_$$7 CDN     VSS     VSS     N      L=0.18U     W=0.83U  
M22     U78_in  u8_D    U75_$$7 VSS     N      L=0.18U     W=0.83U  
M23     U15_S   U15_GB  U77_in  VDD     P      L=0.18U     W=1.38U   PD=.520U
M24     U15_S   U15_G   U77_in  VSS     N      L=0.18U     W=0.42U   PD=.480U
M25     U77_out U15_G   u8_D    VDD     P      L=0.18U     W=0.69U  
M26     U77_out U15_GB  u8_D    VSS     N      L=0.18U     W=0.4U  
M27     U76_out U15_G   U77_in  VDD     P      L=0.189U    W=1.38U  
M28     U76_out U15_GB  U77_in  VSS     N      L=0.18U     W=0.46U  
M29     u9_S    U15_GB  u8_D    VDD     P      L=0.18U     W=0.69U  
M30     u9_S    U15_G   u8_D    VSS     N      L=0.18U     W=0.47U  
M31     U67_drain D       U15_S   VDD     P    L=0.185U    W=1.78U   
+  PS=.520U PD=.520U
M32     VDD     U43_gate U67_drain VDD     P   L=0.185U    W=1.78U   
+  PS=.520U
M33     U66_drain SD      U15_S   VDD     P    L=0.184U    W=1.91U   
+  PS=.520U PD=.520U
M34     VDD     U45_gate U66_drain VDD     P   L=0.184U    W=1.91U   
+  PS=.520U
M35     U68_drain U45_gate VSS     VSS     N   L=0.18U     W=0.69U   
+  PD=.480U
M36     U69_drain U43_gate VSS     VSS     N   L=0.18U     W=.66U   
+  PD=.480U
M37     U15_S   D       U68_drain VSS     N    L=0.18U     W=0.69U   
+  PS=.480U PD=.480U
M38     U15_S   SD      U69_drain VSS     N    L=0.18U     W=.66U   
+  PS=.480U PD=.480U

.ENDS sdcrn4

.SUBCKT sdcrq4 Q  CDN CP D SC SD VDD VSS
M1      U77_out U77_in  VSS     VSS     N   L=0.18U  W=0.82U  
M2      U77_out U77_in  VDD     VDD     P   L=0.18U  W=1.66U  
M3      U15_G   CP      VSS     VSS     N   L=0.18U  W=0.66U  
M4      U15_G   CP      VDD     VDD     P   L=0.184U  W=1.74U  
M5      U15_GB  U15_G   VSS     VSS     N   L=0.18U  W=0.66U  
M6      U15_GB  U15_G   VDD     VDD     P   L=0.184U  W=1.74U  
M7      U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M8      U43_gate U45_gate VDD     VDD     P   L=0.184U  W=1.91U  
M9      U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M10     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M11     U78_out U78_in  VSS     VSS     N   L=0.18U  W=0.83U  
M12     U78_out U78_in  VDD     VDD     P   L=0.185U  W=1.66U  
M13     Q       U78_in  VSS     VSS     N   L=0.18U  W=2.88U  
M14     Q       U78_in  VDD     VDD     P   L=0.184U  W=8.20U  
M15     U76_out CDN     VDD     VDD     P   L=0.18U  W=1.36U  
M16     U76_out U77_out VDD     VDD     P   L=0.18U  W=1.36U  
M17     U76_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.82U  
M18     U76_out U77_out U76_$$7 VSS     N   L=0.18U  W=0.82U  
M19     U78_in  CDN     VDD     VDD     P   L=0.185U  W=1.45U  
M20     U78_in  u8_D    VDD     VDD     P   L=0.18U  W=1.45U  
M21     U75_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.83U  
M22     U78_in  u8_D    U75_$$7 VSS     N   L=0.18U  W=0.83U  
M23     VDD     U45_gate U45_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M24     U67_drain D       U15_S   VDD     P   L=0.18U  W=1.78U   
+  PS=.520U PD=.520U
M25     VDD     U43_gate U67_drain VDD     P   L=0.18U  W=1.78U   
+  PS=.520U
M26     U45_source SD      U15_S   VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M27     U15_S   U15_GB  U77_in  VDD     P   L=0.18U  W=1.38U   PD=.520U
M28     U15_S   U15_G   U77_in  VSS     N   L=0.18U  W=0.42U   PD=.480U
M29     U76_out U15_G   U77_in  VDD     P   L=0.18U  W=1.38U  
M30     U76_out U15_GB  U77_in  VSS     N   L=0.18U  W=0.46U  
M31     U77_out U15_G   u8_D    VDD     P   L=0.18U  W=0.69U  
M32     U77_out U15_GB  u8_D    VSS     N   L=0.18U  W=0.40U  
M33     U78_out U15_GB  u8_D    VDD     P   L=0.18U  W=0.69U  
M34     U78_out U15_G   u8_D    VSS     N   L=0.18U  W=0.47U  
M35     U68_drain U45_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M36     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M37     U15_S   SD      U69_drain VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U
M38     U15_S   D       U68_drain VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U

.ENDS sdcrq4

.SUBCKT sdnfb1 Q QN  CPN D SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.82U  
M2      U35_out U35_in  VDD     VDD     P   L=0.18U  W=1.66U  
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.82U  
M4      U37_out U35_out VDD     VDD     P   L=0.18U  W=1.66U  
M5      u7_G    CPN     VSS     VSS     N   L=0.18U  W=0.66U  
M6      u7_G    CPN     VDD     VDD     P   L=0.184U  W=1.8U  
M7      u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.66U  
M8      u7_GB   u7_G    VDD     VDD     P   L=0.184U  W=1.8U  
M9      U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M10     U43_gate U45_gate VDD     VDD     P   L=0.184U  W=1.91U  
M11     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M12     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M13     u9_S    U36_in  VSS     VSS     N   L=0.18U  W=0.83U  
M14     u9_S    U36_in  VDD     VDD     P   L=0.184U  W=1.88U  
M15     U36_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M16     U36_in  u9_D    VDD     VDD     P   L=0.184U  W=1.88U  
M17     Q       U36_in  VSS     VSS     N   L=0.18U  W=0.75U  
M18     Q       U36_in  VDD     VDD     P   L=0.184U  W=2.05U  
M19     QN      u9_D    VSS     VSS     N   L=0.18U  W=0.75U  
M20     QN      u9_D    VDD     VDD     P   L=0.184U  W=2.05U  
M21     U37_out u7_GB   U35_in  VDD     P   L=0.18U  W=1.25U  
M22     U37_out u7_G    U35_in  VSS     N   L=0.18U  W=0.44U  
M23     U66_source u7_G    U35_in  VDD     P   L=0.18U  W=1.25U   
+  PD=.520U
M24     U66_source u7_GB   U35_in  VSS     N   L=0.18U  W=0.44U   
+  PD=.480U
M25     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.69U  
M26     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M27     U35_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.69U  
M28     U35_out u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  
M29     VDD     U45_gate U45_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M30     U45_source SD      U66_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M31     U67_drain D       U66_source VDD     P   L=0.18U  W=1.78U   
+  PS=.520U PD=.520U
M32     VDD     U43_gate U67_drain VDD     P   L=0.18U  W=1.78U   
+  PS=.520U
M33     U66_source D       U48_source VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M34     U48_source U45_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M35     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M36     U66_source SD      U69_drain VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U

.ENDS sdnfb1

.SUBCKT sdnfb2 Q QN  CPN D SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.82U  
M2      U35_out U35_in  VDD     VDD     P   L=0.18U  W=1.66U  
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.82U  
M4      U37_out U35_out VDD     VDD     P   L=0.18U  W=1.66U  
M5      u7_G    CPN     VSS     VSS     N   L=0.18U  W=0.66U  
M6      u7_G    CPN     VDD     VDD     P   L=0.184U  W=1.8U  
M7      u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.66U  
M8      u7_GB   u7_G    VDD     VDD     P   L=0.184U  W=1.8U  
M9      U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M10     U43_gate U45_gate VDD     VDD     P   L=0.184U  W=1.91U  
M11     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M12     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M13     u9_S    U36_in  VSS     VSS     N   L=0.18U  W=.83U  
M14     u9_S    U36_in  VDD     VDD     P   L=0.184U  W=1.88U  
M15     U36_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M16     U36_in  u9_D    VDD     VDD     P   L=0.184U  W=1.88U  
M17     Q       U36_in  VSS     VSS     N   L=0.18U  W=1.43U  
M18     Q       U36_in  VDD     VDD     P   L=0.182U  W=4.1U  
M19     QN      u9_D    VSS     VSS     N   L=0.18U  W=1.43U  
M20     QN      u9_D    VDD     VDD     P   L=0.184U  W=4.1U  
M21     U37_out u7_GB   U35_in  VDD     P   L=0.18U  W=1.25U  
M22     U37_out u7_G    U35_in  VSS     N   L=0.18U  W=0.44U  
M23     U66_source u7_G    U35_in  VDD     P   L=0.18U  W=1.25U   
+  PD=.520U
M24     U66_source u7_GB   U35_in  VSS     N   L=0.18U  W=0.44U   
+  PD=.480U
M25     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.69U  
M26     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M27     U35_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.69U  
M28     U35_out u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  
M29     VDD     U45_gate U45_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M30     U45_source SD      U66_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M31     U67_drain D       U66_source VDD     P   L=0.18U  W=1.78U   
+  PS=.520U PD=.520U
M32     VDD     U43_gate U67_drain VDD     P   L=0.18U  W=1.78U   
+  PS=.520U
M33     U66_source D       U48_source VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M34     U48_source U45_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M35     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M36     U66_source SD      U69_drain VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U

.ENDS sdnfb2

.SUBCKT sdnfb4 Q QN  CPN D SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.82U  
M2      U35_out U35_in  VDD     VDD     P   L=0.18U  W=1.66U  
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.82U  
M4      U37_out U35_out VDD     VDD     P   L=0.18U  W=1.66U  
M5      u7_G    CPN     VSS     VSS     N   L=0.18U  W=0.66U  
M6      u7_G    CPN     VDD     VDD     P   L=0.184U  W=1.8U  
M7      u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.66U  
M8      u7_GB   u7_G    VDD     VDD     P   L=0.184U  W=1.8U  
M9      U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M10     U43_gate U45_gate VDD     VDD     P   L=0.184U  W=1.91U  
M11     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M12     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M13     u9_S    U36_in  VSS     VSS     N   L=0.18U  W=.83U  
M14     u9_S    U36_in  VDD     VDD     P   L=0.184U  W=1.88U  
M15     U36_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M16     U36_in  u9_D    VDD     VDD     P   L=0.184U  W=1.88U  
M17     Q       U36_in  VSS     VSS     N   L=0.18U  W=2.94U  
M18     Q       U36_in  VDD     VDD     P   L=0.182U  W=8.20U  
M19     QN      u9_D    VSS     VSS     N   L=0.18U  W=2.94U  
M20     QN      u9_D    VDD     VDD     P   L=0.184U  W=8.20U  
M21     U37_out u7_GB   U35_in  VDD     P   L=0.18U  W=1.25U  
M22     U37_out u7_G    U35_in  VSS     N   L=0.18U  W=0.44U  
M23     U66_source u7_G    U35_in  VDD     P   L=0.18U  W=1.25U   
+  PD=.520U
M24     U66_source u7_GB   U35_in  VSS     N   L=0.18U  W=0.44U   
+  PD=.480U
M25     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.69U  
M26     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M27     U35_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.69U  
M28     U35_out u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  
M29     VDD     U45_gate U45_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M30     U45_source SD      U66_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M31     U67_drain D       U66_source VDD     P   L=0.18U  W=1.78U   
+  PS=.520U PD=.520U
M32     VDD     U43_gate U67_drain VDD     P   L=0.18U  W=1.78U   
+  PS=.520U
M33     U66_source D       U48_source VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M34     U48_source U45_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M35     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M36     U66_source SD      U69_drain VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U

.ENDS sdnfb4

.SUBCKT sdnrb4 Q QN  CP D SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.82U  
M2      U35_out U35_in  VDD     VDD     P   L=0.18U  W=1.66U  
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.82U  
M4      U37_out U35_out VDD     VDD     P   L=0.185U  W=1.66U  
M5      u7_GB   CP      VSS     VSS     N   L=0.18U  W=0.66U  
M6      u7_GB   CP      VDD     VDD     P   L=0.184U  W=1.74U  
M7      u7_G    u7_GB   VSS     VSS     N   L=0.18U  W=0.66U  
M8      u7_G    u7_GB   VDD     VDD     P   L=0.184U  W=1.74U  
M9      U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M10     U43_gate U45_gate VDD     VDD     P   L=0.184U  W=1.91U  
M11     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M12     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M13     u9_S    U36_in  VSS     VSS     N   L=0.18U  W=.83U  
M14     u9_S    U36_in  VDD     VDD     P   L=0.184U  W=1.88U  
M15     U36_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M16     U36_in  u9_D    VDD     VDD     P   L=0.184U  W=1.88U  
M17     Q       U36_in  VSS     VSS     N   L=0.18U  W=2.94U  
M18     Q       U36_in  VDD     VDD     P   L=0.182U  W=8.2U  
M19     QN      u9_D    VSS     VSS     N   L=0.18U  W=2.94U  
M20     QN      u9_D    VDD     VDD     P   L=0.182U  W=8.2U  
M21     U37_out u7_GB   U35_in  VDD     P   L=0.18U  W=1.38U  
M22     U37_out u7_G    U35_in  VSS     N   L=0.18U  W=0.46U  
M23     U66_source u7_G    U35_in  VDD     P   L=0.186U  W=1.38U   
+  PD=.520U
M24     U66_source u7_GB   U35_in  VSS     N   L=0.18U  W=0.42U   
+  PD=.480U
M25     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.69U  
M26     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M27     u9_D    u7_GB   U35_out VDD     P   L=0.18U  W=0.69U  
M28     u9_D    u7_G    U35_out VSS     N   L=0.18U  W=0.46U  
M29     VDD     U45_gate U45_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M30     U45_source SD      U66_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M31     U67_drain D       U66_source VDD     P   L=0.185U  W=1.78U   
+  PS=.520U PD=.520U
M32     VDD     U43_gate U67_drain VDD     P   L=0.185U  W=1.78U   
+  PS=.520U
M33     U66_source D       U48_source VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M34     U48_source U45_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M35     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M36     U66_source SD      U69_drain VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U

.ENDS sdnrb4

.SUBCKT sdnrn4 QN  CP D SC SD VDD VSS
M1      u7_S    u7_GB   u7_D    VDD     P   L=.18U      	W=1.38U
M2      u7_S    u7_G    u7_D    VSS     N   L=.18U     		 W=0.46U   
M3      U36_out u7_G    u9_D    VDD     P   L=.18U  		W=0.69U    
M4      U36_out u7_GB   u9_D    VSS     N   L=.18U		  W=0.42U    
M5      U50_drain u7_G    u7_D    VDD     P   L=.186U 		 W=1.38U     
+  PD=.520U
M6      U50_drain u7_GB   u7_D    VSS     N   L=.18U 		 W=0.46U    
+  PD=.480U
M7      u9_D    u7_GB   U37_in  VDD     P   L=.18U 		 W=0.69U    
M8      u9_D    u7_G    U37_in  VSS     N   L=.18U 		 W=0.46U    
M9      VDD     U43_gate U43_source VDD     P   L=.184U  	W=1.78U     
+  PS=.520U
M10     U43_source D       U50_drain VDD     P   L=.184U  	W=1.78U     
+  PS=.520U PD=.520U
M11     VDD     U68_gate U45_source VDD     P   L=.18U  	W=1.91U    
+  PS=.520U
M12     U45_source SD      U50_drain VDD     P   L=.18U 	 W=1.91U     
+  PS=.520U PD=.520U
M13     U36_out U36_in  VSS     VSS     N   L=.18U 		 W=0.83U    
M14     U36_out U36_in  VDD     VDD     P   L=.184U  		W=1.88U    
M15     u7_S    U37_in  VSS     VSS     N   L=.18U 		 W=0.82U    
M16     u7_S    U37_in  VDD     VDD     P   L=.185U  		W=1.66U    
M17     u7_G    u7_GB   VSS     VSS     N   L=.18U  		W=0.66U    
M18     u7_G    u7_GB   VDD     VDD     P   L=.184U  		W=1.74U    
M19     u7_GB   CP      VSS     VSS     N   L=.18U  		W=0.66U   
M20     u7_GB   CP      VDD     VDD     P   L=.18U 		 W=1.74U   
M21     U43_gate U68_gate VSS     VSS     N   L=.18U  		W=0.69U    
M22     U43_gate U68_gate VDD     VDD     P   L=.18U  		W=1.91U   
M23     U68_gate SC      VSS     VSS     N   L=.18U  		W=0.69U    
M24     U68_gate SC      VDD     VDD     P   L=.184U 		 W=1.91U    
M25     U36_in  u9_D    VSS     VSS     N   L=.18U 		 W=0.83U    
M26     U36_in  u9_D    VDD     VDD     P   L=.18U 		 W=1.88U    
M27     U37_in  u7_D    VSS     VSS     N   L=.18U 		 W=0.82U    
M28     U37_in  u7_D    VDD     VDD     P   L=.185U 		 W=1.66U    
M29     QN      u9_D    VSS     VSS     N   L=.184U  		W=2.82U   
M30     QN      u9_D    VDD     VDD     P   L=.182U  		W=8.09U    
M31     U50_drain SD      U50_source VSS     N   L=.18U  	W=0.66U     
+  PS=.480U PD=.480U
M32     U50_source U43_gate VSS     VSS     N   L=.18U  	W=.66U     
+  PD=.480U
M33     U50_drain D       U48_source VSS     N   L=.18U  	W=0.69U     
+  PS=.480U PD=.480U
M34     U48_source U68_gate VSS     VSS     N   L=.18U 		 W=0.69U    
+  PD=.480U

.ENDS sdnrn4

.SUBCKT sdnrq4 Q  CP D SC SD VDD VSS
M1      u7_S    u7_GB   u7_D    VDD     P   L=0.18U  W=1.38U  
M2      u7_S    u7_G    u7_D    VSS     N   L=0.18U  W=0.46U  
M3      U36_out u7_G    u9_D    VDD     P   L=0.18U  W=0.69U  
M4      U36_out u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M5      U50_drain u7_G    u7_D    VDD     P   L=0.186U  W=1.38U   
+  PD=.520U
M6      U50_drain u7_GB   u7_D    VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M7      u9_D    u7_GB   U37_in  VDD     P   L=0.18U  W=0.69U  
M8      u9_D    u7_G    U37_in  VSS     N   L=0.18U  W=0.46U  
M9      VDD     U43_gate U43_source VDD     P   L=0.185U  W=1.78U   
+  PS=.520U
M10     U43_source D       U50_drain VDD     P   L=0.185U  W=1.78U   
+  PS=.520U PD=.520U
M11     VDD     U68_gate U45_source VDD     P   L=0.18U  W=1.91U   
+  PS=.520U
M12     U45_source SD      U50_drain VDD     P   L=0.18U  W=1.91U   
+  PS=.520U PD=.520U
M13     U36_out U36_in  VSS     VSS     N   L=0.18U  W=0.83U  
M14     U36_out U36_in  VDD     VDD     P   L=0.184U  W=1.88U  
M15     u7_S    U37_in  VSS     VSS     N   L=0.18U  W=0.82U  
M16     u7_S    U37_in  VDD     VDD     P   L=0.185U  W=1.66U  
M17     u7_G    u7_GB   VSS     VSS     N   L=0.18U  W=0.66U  
M18     u7_G    u7_GB   VDD     VDD     P   L=0.184U  W=1.74U  
M19     u7_GB   CP      VSS     VSS     N   L=0.18U  W=0.66U  
M20     u7_GB   CP      VDD     VDD     P   L=0.184U  W=1.74U  
M21     U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U  
M22     U43_gate U68_gate VDD     VDD     P   L=0.18U  W=1.91U  
M23     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M24     U68_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M25     Q       U36_in  VSS     VSS     N   L=0.18U  W=2.82U  
M26     Q       U36_in  VDD     VDD     P   L=0.182U  W=8.09U  
M27     U36_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M28     U36_in  u9_D    VDD     VDD     P   L=0.18U  W=1.88U  
M29     U37_in  u7_D    VSS     VSS     N   L=0.18U  W=0.82U  
M30     U37_in  u7_D    VDD     VDD     P   L=0.18U  W=1.66U  
M31     U50_drain SD      U50_source VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U
M32     U50_source U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M33     U50_drain D       U48_source VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M34     U48_source U68_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U

.ENDS sdnrq4

.SUBCKT sdpfb1 Q QN  CPN D SC SD SDN VDD VSS
M1      U37_out U37_in  VSS     VSS     N   L=0.18U  W=0.79U  
M2      U37_out U37_in  VDD     VDD     P   L=0.185U  W=1.83U  
M3      u7_G    CPN     VSS     VSS     N   L=0.18U  W=0.69U  
M4      u7_G    CPN     VDD     VDD     P   L=0.185U  W=1.8U  
M5      u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.69U  
M6      u7_GB   u7_G    VDD     VDD     P   L=0.18U  W=1.8U  
M7      U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M8      U43_gate U45_gate VDD     VDD     P   L=0.18U  W=1.91U  
M9      U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M10     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M11     QN      u9_D    VSS     VSS     N   L=0.18U  W=0.69U  
M12     QN      u9_D    VDD     VDD     P   L=0.185U  W=2.05U  
M13     Q       U74_in1 VSS     VSS     N   L=0.18U  W=0.69U  
M14     Q       U74_in1 VDD     VDD     P   L=0.184U  W=1.969U  
M15     U74_in1 u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M16     U74_in1 u9_D    VDD     VDD     P   L=0.184U  W=1.99U  
M17     U37_in  SDN     VDD     VDD     P   L=0.18U  W=1.38U  
M18     U37_in  U73_in1 VDD     VDD     P   L=0.186U  W=1.38U  
M19     U73_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.83U  
M20     U37_in  U73_in1 U73_$$7 VSS     N   L=0.18U  W=0.83U  
M21     U74_out SDN     VDD     VDD     P   L=0.18U  W=1.38U  
M22     U74_out U74_in1 VDD     VDD     P   L=0.186U  W=1.38U  
M23     U74_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.83U  
M24     U74_out U74_in1 U74_$$7 VSS     N   L=0.18U  W=0.83U  
M25     VDD     U43_gate U43_source VDD     P   L=0.185U  W=1.78U   
+  PS=.520U
M26     U43_source D       U67_source VDD     P   L=0.185U  W=1.78U   
+  PS=.520U PD=.520U
M27     VDD     U45_gate U45_source VDD     P   L=0.18U  W=1.91U   
+  PS=.520U
M28     U45_source SD      U67_source VDD     P   L=0.18U  W=1.91U   
+  PS=.520U PD=.520U
M29     U37_out u7_GB   U73_in1 VDD     P   L=0.18U  W=1.25U  
M30     U37_out u7_G    U73_in1 VSS     N   L=0.18U  W=0.46U  
M31     U67_source u7_G    U73_in1 VDD     P   L=0.187U  W=1.25U   
+  PD=.520U
M32     U67_source u7_GB   U73_in1 VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M33     U74_out u7_G    u9_D    VDD     P   L=0.18U  W=0.83U  
M34     U74_out u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M35     U37_in  u7_GB   u9_D    VDD     P   L=0.18U  W=0.83U  
M36     U37_in  u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  
M37     U67_source D       U48_source VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M38     U48_source U45_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M39     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M40     U67_source SD      U69_drain VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U

.ENDS sdpfb1

.SUBCKT sdpfb2 Q QN  CPN D SC SD SDN VDD VSS
M1      U37_out U37_in  VSS     VSS     N   L=0.18U  W=0.79U    
M2      U37_out U37_in  VDD     VDD     P   L=0.185U  W=1.83U    
M3      u7_G    CPN     VSS     VSS     N   L=0.18U  W=0.69U   
M4      u7_G    CPN     VDD     VDD     P   L=0.185U  W=1.8U    
M5      u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.69U    
M6      u7_GB   u7_G    VDD     VDD     P   L=0.18U  W=1.8U    
M7      U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U    
M8      U43_gate U45_gate VDD     VDD     P   L=0.184U  W=1.91U    
M9      U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U    
M10     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U    
M11     QN      u9_D    VSS     VSS     N   L=0.18U  W=1.38U    
M12     QN      u9_D    VDD     VDD     P   L=0.184U  W=4.1U    
M13     Q       U74_in1 VSS     VSS     N   L=0.18U  W=1.44U    
M14     Q       U74_in1 VDD     VDD     P   L=0.184U  W=4.1U    
M15     U74_in1 u9_D    VSS     VSS     N   L=0.18U  W=0.83U    
M16     U74_in1 u9_D    VDD     VDD     P   L=0.184U  W=1.99U    
M17     U37_in  SDN     VDD     VDD     P   L=0.18U  W=1.38U    
M18     U37_in  U73_in1 VDD     VDD     P   L=0.186U  W=1.38U    
M19     U73_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.79U    
M20     U37_in  U73_in1 U73_$$7 VSS     N   L=0.18U  W=0.79U    
M21     U74_out SDN     VDD     VDD     P   L=0.18U  W=1.38U    
M22     U74_out U74_in1 VDD     VDD     P   L=0.186U  W=1.38U    
M23     U74_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.83U    
M24     U74_out U74_in1 U74_$$7 VSS     N   L=0.18U  W=0.83U    
M25     VDD     U43_gate U43_source VDD     P   L=0.185U  W=1.78U     
+  PS=.520U
M26     U43_source D       U67_source VDD     P   L=0.185U  W=1.78U     
+  PS=.520U PD=.520U
M27     VDD     U45_gate U45_source VDD     P   L=0.184U  W=1.91U     
+  PS=.520U
M28     U45_source SD      U67_source VDD     P   L=0.189U  W=1.91U     
+  PS=.520U PD=.520U
M29     U37_out u7_GB   U73_in1 VDD     P   L=0.18U  W=1.25U    
M30     U37_out u7_G    U73_in1 VSS     N   L=0.18U  W=0.46U    
M31     U67_source u7_G    U73_in1 VDD     P   L=0.187U  W=1.25U     
+  PD=.520U
M32     U67_source u7_GB   U73_in1 VSS     N   L=0.18U  W=0.46U     
+  PD=.480U
M33     U74_out u7_G    u9_D    VDD     P   L=0.18U  W=0.83U    
M34     U74_out u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U    
M35     U37_in  u7_GB   u9_D    VDD     P   L=0.18U  W=0.83U    
M36     U37_in  u7_G    u9_D    VSS     N   L=0.18U  W=0.46U    
M37     U67_source D       U48_source VSS     N   L=0.18U  W=0.69U     
+  PS=.480U PD=.480U
M38     U48_source U45_gate VSS     VSS     N   L=0.18U  W=0.69U     
+  PD=.480U
M39     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U     
+  PD=.480U
M40     U67_source SD      U69_drain VSS     N   L=0.18U  W=0.66U     
+  PS=.480U PD=.480U

.ENDS sdpfb2

.SUBCKT sdpfb4 Q QN  CPN D SC SD SDN VDD VSS
M1      U37_out U37_in  VSS     VSS     N   L=0.18U  W=0.79U    
M2      U37_out U37_in  VDD     VDD     P   L=0.185U  W=1.83U    
M3      u7_G    CPN     VSS     VSS     N   L=0.18U  W=0.69U    
M4      u7_G    CPN     VDD     VDD     P   L=0.185U  W=1.8U    
M5      u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.69U    
M6      u7_GB   u7_G    VDD     VDD     P   L=0.18U  W=1.8U    
M7      U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U    
M8      U43_gate U45_gate VDD     VDD     P   L=0.184U  W=1.91U    
M9      U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U    
M10     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U    
M11     QN      u9_D    VSS     VSS     N   L=0.18U  W=2.94U    
M12     QN      u9_D    VDD     VDD     P   L=0.183U  W=8.2U    
M13     Q       U74_in1 VSS     VSS     N   L=0.18U  W=2.99U    
M14     Q       U74_in1 VDD     VDD     P   L=0.183U  W=8.2U    
M15     U74_in1 u9_D    VSS     VSS     N   L=0.18U  W=0.83U    
M16     U74_in1 u9_D    VDD     VDD     P   L=0.184U  W=1.99U    
M17     U37_in  SDN     VDD     VDD     P   L=0.18U  W=1.38U    
M18     U37_in  U73_in1 VDD     VDD     P   L=0.186U  W=1.38U    
M19     U73_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.79U    
M20     U37_in  U73_in1 U73_$$7 VSS     N   L=0.18U  W=0.79U    
M21     U74_out SDN     VDD     VDD     P   L=0.18U  W=1.38U    
M22     U74_out U74_in1 VDD     VDD     P   L=0.186U  W=1.38U    
M23     U74_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.83U    
M24     U74_out U74_in1 U74_$$7 VSS     N   L=0.18U  W=0.83U    
M25     VDD     U43_gate U43_source VDD     P   L=0.185U  W=1.78U     
+  PS=.520U
M26     U43_source D       U67_source VDD     P   L=0.185U  W=1.78U     
+  PS=.520U PD=.520U
M27     VDD     U45_gate U45_source VDD     P   L=0.184U  W=1.91U     
+  PS=.520U
M28     U45_source SD      U67_source VDD     P   L=0.189U  W=1.91U     
+  PS=.520U PD=.520U
M29     U37_out u7_GB   U73_in1 VDD     P   L=0.18U  W=1.25U    
M30     U37_out u7_G    U73_in1 VSS     N   L=0.18U  W=0.46U    
M31     U67_source u7_G    U73_in1 VDD     P   L=0.187U  W=1.25U     
+  
M32     U67_source u7_GB   U73_in1 VSS     N   L=0.18U  W=0.46U     
+  PD=.480U
M33     U74_out u7_G    u9_D    VDD     P   L=0.18U  W=0.83U    
M34     U74_out u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U    
M35     U37_in  u7_GB   u9_D    VDD     P   L=0.18U  W=0.83U    
M36     U37_in  u7_G    u9_D    VSS     N   L=0.18U  W=0.46U    
M37     U67_source D       U48_source VSS     N   L=0.18U  W=0.69U     
+  PS=.480U PD=.480U
M38     U48_source U45_gate VSS     VSS     N   L=0.18U  W=0.69U     
+  PD=.480U
M39     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U     
+  PD=.480U
M40     U67_source SD      U69_drain VSS     N   L=0.18U  W=0.66U     
+  PS=.480U PD=.480U

.ENDS sdpfb4

.SUBCKT sdprb4 Q QN  CP D SC SD SDN VDD VSS
M1      U37_out U37_in  VSS     VSS     N   L=0.18U  W=0.82U  
M2      U37_out U37_in  VDD     VDD     P   L=0.185U  W=1.8U  
M3      u7_GB   CP      VSS     VSS     N   L=0.18U  W=0.66U  
M4      u7_GB   CP      VDD     VDD     P   L=0.185U  W=1.74U  
M5      u7_G    u7_GB   VSS     VSS     N   L=0.18U  W=0.66U  
M6      u7_G    u7_GB   VDD     VDD     P   L=0.18U  W=1.74U  
M7      U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M8      U43_gate U45_gate VDD     VDD     P   L=0.18U  W=1.91U  
M9      U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M10     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M11     Q       U74_in1 VSS     VSS     N   L=0.18U  W=2.94U  
M12     Q       U74_in1 VDD     VDD     P   L=0.182U  W=8.2U  
M13     U74_in1 u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M14     U74_in1 u9_D    VDD     VDD     P   L=0.18U  W=1.94U  
M15     QN      u9_D    VSS     VSS     N   L=0.18U  W=2.94U  
M16     QN      u9_D    VDD     VDD     P   L=0.18225U  W=8.2U  
M17     U37_in  SDN     VDD     VDD     P   L=0.18U  W=1.38U  
M18     U37_in  U73_in1 VDD     VDD     P   L=0.185U  W=1.38U  
M19     U73_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.82U  
M20     U37_in  U73_in1 U73_$$7 VSS     N   L=0.18U  W=0.82U  
M21     U74_out SDN     VDD     VDD     P   L=0.18U  W=1.38U  
M22     U74_out U74_in1 VDD     VDD     P   L=0.185U  W=1.38U  
M23     U74_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.83U  
M24     U74_out U74_in1 U74_$$7 VSS     N   L=0.18U  W=0.83U  
M25     VDD     U43_gate U43_source VDD     P   L=0.18U  W=1.78U   
+  PS=.520U
M26     VDD     U45_gate U45_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M27     U45_source SD      U66_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M28     U43_source D       U66_source VDD     P   L=0.18U  W=1.78U   
+  PS=.520U PD=.520U
M29     U37_out u7_GB   U73_in1 VDD     P   L=0.18U  W=1.11U  
M30     U37_out u7_G    U73_in1 VSS     N   L=0.18U  W=0.46U  
M31     U66_source u7_G    U73_in1 VDD     P   L=0.18U  W=1.11U   
+  PD=.520U
M32     U66_source u7_GB   U73_in1 VSS     N   L=0.18U  W=0.42U   
+  PD=.480U
M33     U74_out u7_G    u9_D    VDD     P   L=0.18U  W=0.78U  
M34     U74_out u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M35     U37_in  u7_GB   u9_D    VDD     P   L=0.18U  W=0.78U  
M36     U37_in  u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  
M37     U66_source D       U48_source VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M38     U48_source U45_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M39     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U   
+  PD=.480U
M40     U66_source SD      U69_drain VSS     N   L=0.18U  W=0.66U   
+  PS=.480U PD=.480U

.ENDS sdprb4

.SUBCKT secfq1 Q  CDN CPN D ENN SC SD VDD VSS
M1      U22_out QmN     VSS     VSS     N   L=.180U  W=0.61U  
M2      U22_out QmN     VDD     VDD     P   L=.180U  W=1.21U  
M3      U125_out CPN     VSS     VSS     N   L=.180U  W=0.83U  
M4      U125_out CPN     VDD     VDD     P   L=.184U  W=1.932U  
M5      U118_gate ENN     VSS     VSS     N   L=.180U  W=0.72U  
M6      U118_gate ENN     VDD     VDD     P   L=.1840U  W=1.68U  
M7      U120_gate SC      VSS     VSS     N   L=.180U  W=0.83U  
M8      U120_gate SC      VDD     VDD     P   L=.183U  W=2.08U  
M9      U108_gate U120_gate VSS     VSS     N   L=.180U  W=0.71U  
M10     U108_gate U120_gate VDD     VDD     P   L=.183U  W=2.08U  
M11     u7_GB   U125_out VSS     VSS     N   L=.180U  W=0.84U  
M12     u7_GB   U125_out VDD     VDD     P   L=.184U  W=1.92U  
M13     U119_gate U130_out VSS     VSS     N   L=.180U  W=.83U  
M14     U119_gate U130_out VDD     VDD     P   L=.180U  W=1.66U  
M15     Q       U130_out VSS     VSS     N   L=.180U  W=0.69U  
M16     Q       U130_out VDD     VDD     P   L=.180U  W=2.05U  
M17     U119_drain U119_gate DmN     VDD     P   L=.185U  W=1.45U   
+  PS=.750U PD=.750U
M18     U115_drain ENN     U115_source VDD     P   L=.180U  W=1.74U   
+  PS=.750U PD=.750U
M19     U115_source D       DmN     VDD     P   L=.184U  W=1.74U   
+  PS=.750U PD=.750U
M20     VDD     U108_gate U115_drain VDD     P   L=.180U  W=1.40U   
+  PS=.750U
M21     VDD     U108_gate U117_source VDD     P   L=.185U  W=1.45U   
+  PS=.750U
M22     U117_source U118_gate U119_drain VDD     P   L=.180U  W=1.45U  
+   PS=.750U PD=.750U
M23     U102_drain SD      DmN     VDD     P   L=.180U  W=1.3U   
+  PS=.750U PD=.750U
M24     VDD     U120_gate U102_drain VDD     P   L=.180U  W=1.44U   
+  PS=.750U
M25     U120_drain U120_gate VSS     VSS     N   L=.180U  W=0.83U   
+  PD=.500U
M26     U121_drain ENN     U120_drain VSS     N   L=.180U  W=0.76U   
+  PS=.500U PD=.500U
M27     DmN     U119_gate U121_drain VSS     N   L=.180U  W=0.83U   
+  PS=.500U PD=.500U
M28     U104_drain U120_gate VSS     VSS     N   L=.180U  W=.69U   
+  PD=.500U
M29     DmN     SD      U105_source VSS     N   L=.180U  W=0.71U   
+  PS=.500U PD=.500U
M30     U105_source U108_gate VSS     VSS     N   L=.180U  W=0.71U   
+  PD=.500U
M31     DmN     D       U106_source VSS     N   L=.180U  W=.69U   
+  PS=.500U PD=.500U
M32     U106_source U118_gate U104_drain VSS     N   L=.180U  W=.69U  
+   PS=.500U PD=.500U
M33     u7_S    u7_GB   QmN     VDD     P   L=.185U  W=1.36U  
M34     u7_S    U125_out QmN     VSS     N   L=.180U  W=0.80U  
M35     DmN     U125_out QmN     VDD     P   L=.180U  W=1.36U   
+  PD=.750U
M36     DmN     u7_GB   QmN     VSS     N   L=.180U  W=0.68U   PD=.500U
M37     U22_out u7_GB   U130_in1 VDD     P   L=.186U  W=1.21U  
M38     U22_out U125_out U130_in1 VSS     N   L=.180U  W=0.60U  
M39     U119_gate U125_out U130_in1 VDD     P   L=.186U  W=1.21U  
M40     U119_gate u7_GB   U130_in1 VSS     N   L=.180U  W=0.60U  
M41     U130_out CDN     VDD     VDD     P   L=.186U  W=1.811U  
M42     U130_out U130_in1 VDD     VDD     P   L=.185U  W=1.807U  
M43     U130_$$7 CDN     VSS     VSS     N   L=.180U  W=1.09U  
M44     U130_out U130_in1 U130_$$7 VSS     N   L=.180U  W=1.09U  
M45     u7_S    CDN     VDD     VDD     P   L=.180U  W=1.47U  
M46     u7_S    U22_out VDD     VDD     P   L=.180U  W=1.47U  
M47     U129_$$7 CDN     VSS     VSS     N   L=.180U  W=0.84U  
M48     u7_S    U22_out U129_$$7 VSS     N   L=.180U  W=0.84U  

.ENDS secfq1

.SUBCKT secfq2 Q  CDN CPN D ENN SC SD VDD VSS
M1      U22_out QmN     VSS     VSS     N   L=.180U  W=0.73U  
M2      U22_out QmN     VDD     VDD     P   L=.180U  W=1.21U  
M3      U125_out CPN     VSS     VSS     N   L=.180U  W=0.83U  
M4      U125_out CPN     VDD     VDD     P   L=.183U  W=1.99U  
M5      U118_gate ENN     VSS     VSS     N   L=.180U  W=0.64U  
M6      U118_gate ENN     VDD     VDD     P   L=.184U  W=1.68U  
M7      U120_gate SC      VSS     VSS     N   L=.180U  W=0.73U  
M8      U120_gate SC      VDD     VDD     P   L=.184U  W=1.56U  
M9      U108_gate U120_gate VSS     VSS     N   L=.180U  W=0.81U  
M10     U108_gate U120_gate VDD     VDD     P   L=.184U  W=1.56U  
M11     u7_GB   U125_out VSS     VSS     N   L=.180U  W=0.84U  
M12     u7_GB   U125_out VDD     VDD     P   L=.180U  W=1.92U  
M13     U119_gate U130_out VSS     VSS     N   L=.180U  W=0.66U  
M14     U119_gate U130_out VDD     VDD     P   L=.180U  W=1.66U  
M15     Q       U130_out VSS     VSS     N   L=.180U  W=1.41U  
M16     Q       U130_out VDD     VDD     P   L=.182U  W=4.04U  
M17     U119_drain U119_gate DmN     VDD     P   L=.185U  W=1.45U   
+  PS=.750U PD=.750U
M18     U115_drain ENN     U115_source VDD     P   L=.180U  W=1.74U   
+  PS=.750U PD=.750U
M19     U115_source D       DmN     VDD     P   L=.184U  W=1.74U   
+  PS=.750U PD=.750U
M20     VDD     U108_gate U115_drain VDD     P   L=.180U  W=1.40U   
+  PS=.750U
M21     VDD     U108_gate U117_source VDD     P   L=.185U  W=1.45U   
+  PS=.750U
M22     U117_source U118_gate U119_drain VDD     P   L=.180U  W=1.45U  
+   PS=.750U PD=.750U
M23     U102_drain SD      DmN     VDD     P   L=.180U  W=1.23U   
+  PS=.750U PD=.750U
M24     VDD     U120_gate U102_drain VDD     P   L=.180U  W=1.44U   
+  PS=.750U
M25     U120_drain U120_gate VSS     VSS     N   L=.180U  W=0.60U   
+  PD=.500U
M26     U121_drain ENN     U120_drain VSS     N   L=.180U  W=0.75U   
+  PS=.500U PD=.500U
M27     DmN     U119_gate U121_drain VSS     N   L=.180U  W=0.83U   
+  PS=.500U PD=.500U
M28     U104_drain U120_gate VSS     VSS     N   L=.180U  W=.69U   
+  PD=.500U
M29     DmN     SD      U105_source VSS     N   L=.180U  W=0.71U   
+  PS=.500U PD=.500U
M30     U105_source U108_gate VSS     VSS     N   L=.180U  W=0.71U   
+  PD=.500U
M31     DmN     D       U106_source VSS     N   L=.180U  W=.69U   
+  PS=.500U PD=.500U
M32     U106_source U118_gate U104_drain VSS     N   L=.180U  W=.69U  
+   PS=.500U PD=.500U
M33     u7_S    u7_GB   QmN     VDD     P   L=.185U  W=1.36U  
M34     u7_S    U125_out QmN     VSS     N   L=.180U  W=0.94U  
M35     DmN     U125_out QmN     VDD     P   L=.180U  W=1.36U   
+  PD=.750U
M36     DmN     u7_GB   QmN     VSS     N   L=.180U  W=0.94U   PD=.500U
M37     U22_out u7_GB   U130_in1 VDD     P   L=.186U  W=1.21U  
M38     U22_out U125_out U130_in1 VSS     N   L=.180U  W=0.60U  
M39     U119_gate U125_out U130_in1 VDD     P   L=.186U  W=1.21U  
M40     U119_gate u7_GB   U130_in1 VSS     N   L=.180U  W=0.60U
M41     U130_out CDN     VDD     VDD     P   L=.180U  W=1.72U  
M42     U130_out U130_in1 VDD     VDD     P   L=.180U  W=1.72U  
M43     U130_$$7 CDN     VSS     VSS     N   L=.180U  W=1.09U  
M44     U130_out U130_in1 U130_$$7 VSS     N   L=.180U  W=1.09U  
M45     u7_S    CDN     VDD     VDD     P   L=.180U  W=1.47U  
M46     u7_S    U22_out VDD     VDD     P   L=.180U  W=1.47U  
M47     U129_$$7 CDN     VSS     VSS     N   L=.180U  W=0.94U  
M48     u7_S    U22_out U129_$$7 VSS     N   L=.180U  W=0.94U  

.ENDS secfq2

.SUBCKT secfq4 Q  CDN CPN D ENN SC SD VDD VSS
M1      U22_out QmN     VSS     VSS     N   L=.180U  W=0.61U  
M2      U22_out QmN     VDD     VDD     P   L=.180U  W=1.21U  
M3      U125_out CPN     VSS     VSS     N   L=.180U  W=0.83U  
M4      U125_out CPN     VDD     VDD     P   L=.183U  W=1.99U  
M5      U118_gate ENN     VSS     VSS     N   L=.180U  W=0.72U  
M6      U118_gate ENN     VDD     VDD     P   L=.184U  W=1.68U  
M7      U120_gate SC      VSS     VSS     N   L=.180U  W=0.83U  
M8      U120_gate SC      VDD     VDD     P   L=.183U  W=2.08U  
M9      U108_gate U120_gate VSS     VSS     N   L=.180U  W=0.71U  
M10     U108_gate U120_gate VDD     VDD     P   L=.183U  W=2.08U  
M11     u7_GB   U125_out VSS     VSS     N   L=.180U  W=0.84U  
M12     u7_GB   U125_out VDD     VDD     P   L=.182U  W=1.92U  
M13     U119_gate U130_out VSS     VSS     N   L=.180U  W=.83U  
M14     U119_gate U130_out VDD     VDD     P   L=.180U  W=1.66U  
M15     Q       U130_out VSS     VSS     N   L=.180U  W=2.95U  
M16     Q       U130_out VDD     VDD     P   L=.182U  W=8.21U  
M17     U119_drain U119_gate DmN     VDD     P   L=.185U  W=1.45U   
+  PS=.750U PD=.750U
M18     U115_drain ENN     U115_source VDD     P   L=.180U  W=1.74U   
+  PS=.750U PD=.750U
M19     U115_source D       DmN     VDD     P   L=.1840U  W=1.74U   
+  PS=.750U PD=.750U
M20     VDD     U108_gate U115_drain VDD     P   L=.180U  W=1.40U   
+  PS=.750U
M21     VDD     U108_gate U117_source VDD     P   L=.185U  W=1.45U   
+  PS=.750U
M22     U117_source U118_gate U119_drain VDD     P   L=.180U  W=1.45U  
+   PS=.750U PD=.750U
M23     U102_drain SD      DmN     VDD     P   L=.180U  W=1.30U   
+  PS=.750U PD=.750U
M24     VDD     U120_gate U102_drain VDD     P   L=.180U  W=1.44U   
+  PS=.750U
M25     U120_drain U120_gate VSS     VSS     N   L=.180U  W=0.83U   
+  PD=.500U
M26     U121_drain ENN     U120_drain VSS     N   L=.180U  W=0.76U   
+  PS=.500U PD=.500U
M27     DmN     U119_gate U121_drain VSS     N   L=.180U  W=0.83U   
+  PS=.500U PD=.500U
M28     U104_drain U120_gate VSS     VSS     N   L=.180U  W=.69U   
+  PD=.500U
M29     DmN     SD      U105_source VSS     N   L=.180U  W=0.71U   
+  PS=.500U PD=.500U
M30     U105_source U108_gate VSS     VSS     N   L=.180U  W=0.71U   
+  PD=.500U
M31     DmN     D       U106_source VSS     N   L=.180U  W=.69U   
+  PS=.500U PD=.500U
M32     U106_source U118_gate U104_drain VSS     N   L=.180U  W=.69U  
+   PS=.500U PD=.500U
M33     u7_S    u7_GB   QmN     VDD     P   L=.185U  W=1.36U  
M34     u7_S    U125_out QmN     VSS     N   L=.180U  W=0.80U  
M35     DmN     U125_out QmN     VDD     P   L=.180U  W=1.36U   
+  PD=.750U
M36     DmN     u7_GB   QmN     VSS     N   L=.180U  W=0.68U   PD=.500U
M37     U22_out u7_GB   U130_in1 VDD     P   L=.186U  W=1.21U  
M38     U22_out U125_out U130_in1 VSS     N   L=.180U  W=0.60U  
M39     U119_gate U125_out U130_in1 VDD     P   L=.186U  W=1.21U  
M40     U119_gate u7_GB   U130_in1 VSS     N   L=.180U  W=0.60U  
M41     U130_out CDN     VDD     VDD     P   L=.185U  W=1.815U  
M42     U130_out U130_in1 VDD     VDD     P   L=.185U  W=1.815U  
M43     U130_$$7 CDN     VSS     VSS     N   L=.180U  W=1.09U  
M44     U130_out U130_in1 U130_$$7 VSS     N   L=.180U  W=1.09U  
M45     u7_S    CDN     VDD     VDD     P   L=.180U  W=1.47U  
M46     u7_S    U22_out VDD     VDD     P   L=.180U  W=1.47U  
M47     U129_$$7 CDN     VSS     VSS     N   L=.180U  W=0.84U  
M48     u7_S    U22_out U129_$$7 VSS     N   L=.180U  W=0.84U  

.ENDS secfq4

.SUBCKT secrq4 Q  CDN CP D ENN SC SD VDD VSS
M1      U22_out QmN     VSS     VSS     N   L=.18U  W=0.64U  
M2      U22_out QmN     VDD     VDD     P   L=.186U  W=1.27U  
M3      U125_out CP      VSS     VSS     N   L=.18U  W=0.69U  
M4      U125_out CP      VDD     VDD     P   L=.184U  W=1.78U  
M5      U118_gate ENN     VSS     VSS     N   L=.18U  W=0.72U  
M6      U118_gate ENN     VDD     VDD     P   L=.185U  W=1.68U  
M7      U120_gate SC      VSS     VSS     N   L=.18U  W=0.83U  
M8      U120_gate SC      VDD     VDD     P   L=.185U  W=2.08U  
M9      U108_gate U120_gate VSS     VSS     N   L=.18U  W=0.71U  
M10     U108_gate U120_gate VDD     VDD     P   L=.184U  W=2.08U  
M11     u7_G    U125_out VSS     VSS     N   L=.18U  W=0.69U  
M12     u7_G    U125_out VDD     VDD     P   L=.185U  W=1.71U  
M13     U122_gate U130_out VSS     VSS     N   L=.18U  W=0.83U  
M14     U122_gate U130_out VDD     VDD     P   L=.18U  W=1.66U  
M15     Q       U130_out VSS     VSS     N   L=.183U  W=2.95U  
M16     Q       U130_out VDD     VDD     P   L=.182U  W=8.2U  
M17     U120_drain U120_gate VSS     VSS     N   L=.180U  W=0.83U   
+  PD=.500U
M18     U121_drain ENN     U120_drain VSS     N   L=.18U  W=0.76U   
+  PS=.500U PD=.500U
M19     DmN     U122_gate U121_drain VSS     N   L=.18U  W=0.83U   
+  PS=.500U PD=.500U
M20     U104_drain U120_gate VSS     VSS     N   L=.18U  W=0.69U   
+  PD=.500U
M21     U103_drain U108_gate VSS     VSS     N   L=.18U  W=0.71U   
+  PD=.500U
M22     DmN     SD      U103_drain VSS     N   L=.18U  W=0.71U   
+  PS=.500U PD=.500U
M23     U116_drain U118_gate U104_drain VSS     N   L=.18U  W=0.69U   
+  PS=.500U PD=.500U
M24     DmN     D       U116_drain VSS     N   L=.18U  W=0.69U   
+  PS=.500U PD=.500U
M25     U115_drain ENN     U115_source VDD     P   L=.184U  W=1.74U   
+  PS=.750U PD=.750U
M26     U115_source D       DmN     VDD     P   L=.184U  W=1.74U   
+  PS=.750U PD=.750U
M27     VDD     U108_gate U115_drain VDD     P   L=.18U  W=1.4U   
+  PS=.750U
M28     VDD     U108_gate U117_source VDD     P   L=.185U  W=1.45U   
+  PS=.750U
M29     U117_source U118_gate U118_source VDD     P   L=.185U  W=1.45U 
+    PS=.750U PD=.750U
M30     U118_source U122_gate DmN     VDD     P   L=.18U  W=1.45U   
+  PS=.750U PD=.750U
M31     U102_drain SD      DmN     VDD     P   L=.18U  W=1.3U   
+  PS=.750U PD=.750U
M32     VDD     U120_gate U102_drain VDD     P   L=.185U  W=1.44U   
+  PS=.750U
M33     u7_S    U125_out QmN     VDD     P   L=.18U  W=1.08U  
M34     u7_S    u7_G    QmN     VSS     N   L=.18U  W=0.83U  
M35     DmN     u7_G    QmN     VDD     P   L=.187U  W=1.08U   
+  PD=.750U
M36     DmN     U125_out QmN     VSS     N   L=.18U  W=0.83U   
+  PD=.500U
M37     U22_out U125_out U130_in1 VDD     P   L=.180U  W=1.08U  
M38     U22_out u7_G    U130_in1 VSS     N   L=.180U  W=0.64U  
M39     U122_gate u7_G    U130_in1 VDD     P   L=.187U  W=1.08U  
M40     U122_gate U125_out U130_in1 VSS     N   L=.18U  W=0.69U  
M41     U130_out CDN     VDD     VDD     P   L=.186U  W=1.25U  
M42     U130_out U130_in1 VDD     VDD     P   L=.18U  W=1.63U  
M43     U130_$$7 CDN     VSS     VSS     N   L=.18U  W=0.93U  
M44     U130_out U130_in1 U130_$$7 VSS     N   L=.18U  W=0.93U  
M45     u7_S    CDN     VDD     VDD     P   L=.185U  W=1.45U  
M46     u7_S    U22_out VDD     VDD     P   L=.185U  W=1.45U  
M47     U129_$$7 CDN     VSS     VSS     N   L=.18U  W=0.83U  
M48     u7_S    U22_out U129_$$7 VSS     N   L=.18U  W=0.83U  

.ENDS secrq4

.SUBCKT senrb1 Q QN  D SD CP ENN SC VDD VSS
M1      U128_out U128_in VSS     VSS     N   L=.18U      W=0.83U
M2      U128_out U128_in VDD     VDD     P   L=.184U      W=1.73U
M3      U128_in QmN     VSS     VSS     N   L=.18U     W=0.83U
M4      U128_in QmN     VDD     VDD     P   L=.184U     W=1.73U
M5      U125_out CP      VSS     VSS     N   L=.18U      W=0.69U
M6      U125_out CP      VDD     VDD     P   L=.184U     W=1.77U
M7      U118_gate ENN     VSS     VSS     N   L=.18U     W=0.72U
M8      U118_gate ENN     VDD     VDD     P   L=.18U     W=1.68U
M9      U120_gate SC      VSS     VSS     N   L=.18U     W=0.69U
M10     U120_gate SC      VDD     VDD     P   L=.184U      W=1.76U
M11     U108_gate U120_gate VSS     VSS     N   L=.18U     W=0.69U
M12     U108_gate U120_gate VDD     VDD     P   L=.18U     W=1.76U
M13     U15_GB  U125_out VSS     VSS     N   L=.18U     W=0.68U
M14     U15_GB  U125_out VDD     VDD     P   L=.18U     W=1.25U
M15     U122_gate U23_in  VSS     VSS     N   L=.18U     W=0.83U
M16     U122_gate U23_in  VDD     VDD     P   L=.184U      W=2.22U
M17     U23_in  Qsl     VSS     VSS     N   L=.18U      W=0.83U
M18     U23_in  Qsl     VDD     VDD     P   L=.184U      W=2.22U
M19     Q       U23_in  VSS     VSS     N   L=.18U      W=0.69U
M20     Q       U23_in  VDD     VDD     P   L=.184U     W=2.05U
M21     QN      Qsl     VSS     VSS     N   L=.18U      W=0.69U
M22     QN      Qsl     VDD     VDD     P   L=.184U      W=2.05U
M23     U115_drain ENN     U115_source VDD     P   L=.185U      W=1.4U
+  PS=.750U PD=.750U
M24     U115_source D       DmN     VDD     P   L=.185U      W=1.4U
+  PS=.750U PD=.750U
M25     VDD     U108_gate U115_drain VDD     P   L=.185U      W=1.4U
+  PS=.750U
M26     VDD     U108_gate U117_source VDD     P   L=.185U      W=1.4U
+  PS=.750U
M27     U117_source U118_gate U118_source VDD     P   L=.185U   W=1.4U
+    PS=.750U PD=.750U
M28     U118_source U122_gate DmN     VDD     P   L=.18U      W=1.57U
+  PS=.750U PD=.750U
M29     VDD     U120_gate U109_source VDD     P   L=.18U      W=1.44U
+  PS=.750U
M30     U109_source SD      DmN     VDD     P   L=.18U       W=1.44U
+  PS=.750U PD=.750U
M31     U121_drain ENN     U121_source VSS     N   L=.18U      W=0.72U
+  PS=.500U PD=.500U
M32     DmN     U122_gate U121_drain VSS     N   L=.18U      W=0.83U
+  PS=.500U PD=.500U
M33     U121_source U120_gate VSS     VSS     N   L=.18U      W=0.69U
+  PD=.500U
M34     DmN     D       U106_source VSS     N   L=.18U      W=0.69U
+  PS=.500U PD=.500U
M35     U104_drain U120_gate VSS     VSS     N   L=.18U      W=0.69U
+  PD=.500U
M36     U106_source U118_gate U104_drain VSS     N   L=.18U     W=0.69U
+   PS=.500U PD=.500U
M37     U103_drain U108_gate VSS     VSS     N   L=.18U      W=0.71U
+  PD=.500U
M38     DmN     SD      U103_drain VSS     N   L=.18U      W=0.71U
+  PS=.500U PD=.500U
M39     DmN     U15_GB  QmN     VDD     P   L=.187U      W=1.08U
+  PD=.750U
M40     DmN     U125_out QmN     VSS     N   L=.18U      W=1.04U
+  PD=.500U
M41     U128_out U125_out QmN     VDD     P   L=.187U     W=1.08U
M42     U128_out U15_GB  QmN     VSS     N   L=.18U      W=0.83U
M43     U128_in U125_out Qsl     VDD     P   L=.18U     W=1.08U
M44     U128_in U15_GB  Qsl     VSS     N   L=.18U     W=0.69U
M45     U122_gate U15_GB  Qsl     VDD     P   L=.18U     W=1.08U
M46     U122_gate U125_out Qsl     VSS     N   L=.18U    W=0.69U

.ENDS senrb1

.SUBCKT senrb2 Q QN  D SD CP ENN SC VDD VSS
M1      U128_out U128_in VSS     VSS     N   L=.18U      W=0.83U
M2      U128_out U128_in VDD     VDD     P   L=.184U      W=1.73U
M3      U128_in QmN     VSS     VSS     N   L=.18U     W=0.83U
M4      U128_in QmN     VDD     VDD     P   L=.184U     W=1.73U
M5      U125_out CP      VSS     VSS     N   L=.18U      W=0.69U
M6      U125_out CP      VDD     VDD     P   L=.184U     W=1.77U
M7      U118_gate ENN     VSS     VSS     N   L=.18U     W=0.72U
M8      U118_gate ENN     VDD     VDD     P   L=.18U     W=1.68U
M9      U120_gate SC      VSS     VSS     N   L=.18U     W=0.69U
M10     U120_gate SC      VDD     VDD     P   L=.184U      W=1.76U
M11     U108_gate U120_gate VSS     VSS     N   L=.18U     W=0.69U
M12     U108_gate U120_gate VDD     VDD     P   L=.18U     W=1.76U
M13     U15_GB  U125_out VSS     VSS     N   L=.18U     W=0.68U
M14     U15_GB  U125_out VDD     VDD     P   L=.18U     W=1.25U
M15     U122_gate U23_in  VSS     VSS     N   L=.18U     W=0.83U
M16     U122_gate U23_in  VDD     VDD     P   L=.184U      W=2.22U
M17     U23_in  Qsl     VSS     VSS     N   L=.18U      W=0.83U
M18     U23_in  Qsl     VDD     VDD     P   L=.184U      W=2.22U
M19     Q       U23_in  VSS     VSS     N   L=.18U      W=1.41U
M20     Q       U23_in  VDD     VDD     P   L=.182U     W=4.1U
M21     QN      Qsl     VSS     VSS     N   L=.18U      W=1.41U
M22     QN      Qsl     VDD     VDD     P   L=.182U      W=4.1U
M23     U115_drain ENN     U115_source VDD     P   L=.185U      W=1.4U
+  PS=.750U PD=.750U
M24     U115_source D       DmN     VDD     P   L=.185U      W=1.4U
+  PS=.750U PD=.750U
M25     VDD     U108_gate U115_drain VDD     P   L=.185U      W=1.4U
+  PS=.750U
M26     VDD     U108_gate U117_source VDD     P   L=.185U      W=1.4U
+  PS=.750U
M27     U117_source U118_gate U118_source VDD     P   L=.185U   W=1.4U
+    PS=.750U PD=.750U
M28     U118_source U122_gate DmN     VDD     P   L=.18U      W=1.57U
+  PS=.750U PD=.750U
M29     VDD     U120_gate U109_source VDD     P   L=.18U      W=1.44U
+  PS=.750U
M30     U109_source SD      DmN     VDD     P   L=.18U       W=1.44U
+  PS=.750U PD=.750U
M31     U121_drain ENN     U121_source VSS     N   L=.18U      W=0.72U
+  PS=.500U PD=.500U
M32     DmN     U122_gate U121_drain VSS     N   L=.18U      W=0.83U
+  PS=.500U PD=.500U
M33     U121_source U120_gate VSS     VSS     N   L=.18U      W=0.69U
+  PD=.500U
M34     DmN     D       U106_source VSS     N   L=.18U      W=0.69U
+  PS=.500U PD=.500U
M35     U104_drain U120_gate VSS     VSS     N   L=.18U      W=0.69U
+  PD=.500U
M36     U106_source U118_gate U104_drain VSS     N   L=.18U     W=0.69U
+   PS=.500U PD=.500U
M37     U103_drain U108_gate VSS     VSS     N   L=.18U      W=0.71U
+  PD=.500U
M38     DmN     SD      U103_drain VSS     N   L=.18U      W=0.71U
+  PS=.500U PD=.500U
M39     DmN     U15_GB  QmN     VDD     P   L=.18U      W=1.08U
+  PD=.750U
M40     DmN     U125_out QmN     VSS     N   L=.18U      W=1.04U
+  PD=.500U
M41     U128_out U125_out QmN     VDD     P   L=.187U     W=1.08U
M42     U128_out U15_GB  QmN     VSS     N   L=.18U      W=0.83U
M43     U128_in U125_out Qsl     VDD     P   L=.18U     W=1.08U
M44     U128_in U15_GB  Qsl     VSS     N   L=.18U     W=0.69U
M45     U122_gate U15_GB  Qsl     VDD     P   L=.18U     W=1.08U
M46     U122_gate U125_out Qsl     VSS     N   L=.18U    W=0.69U

.ENDS senrb2

.SUBCKT senrb4 Q QN  D SD CP ENN SC VDD VSS
M1      U128_out U128_in VSS     VSS     N   L=.18U      W=0.83U
M2      U128_out U128_in VDD     VDD     P   L=.184U      W=1.73U
M3      U128_in QmN     VSS     VSS     N   L=.18U     W=0.83U
M4      U128_in QmN     VDD     VDD     P   L=.184U     W=1.73U
M5      U125_out CP      VSS     VSS     N   L=.18U      W=0.69U
M6      U125_out CP      VDD     VDD     P   L=.184U     W=1.77U
M7      U118_gate ENN     VSS     VSS     N   L=.18U     W=0.72U
M8      U118_gate ENN     VDD     VDD     P   L=.18U     W=1.68U
M9      U120_gate SC      VSS     VSS     N   L=.18U     W=0.69U
M10     U120_gate SC      VDD     VDD     P   L=.184U      W=1.76U
M11     U108_gate U120_gate VSS     VSS     N   L=.18U     W=0.69U
M12     U108_gate U120_gate VDD     VDD     P   L=.18U     W=1.76U
M13     U15_GB  U125_out VSS     VSS     N   L=.18U     W=0.68U
M14     U15_GB  U125_out VDD     VDD     P   L=.18U     W=1.25U
M15     U122_gate U23_in  VSS     VSS     N   L=.18U     W=0.83U
M16     U122_gate U23_in  VDD     VDD     P   L=.184U      W=2.22U
M17     U23_in  Qsl     VSS     VSS     N   L=.18U      W=0.83U
M18     U23_in  Qsl     VDD     VDD     P   L=.183U      W=2.22U
M19     Q       U23_in  VSS     VSS     N   L=.18U      W=2.88U
M20     Q       U23_in  VDD     VDD     P   L=.182U     W=8.2U
M21     QN      Qsl     VSS     VSS     N   L=.18U      W=2.88U
M22     QN      Qsl     VDD     VDD     P   L=.182U      W=8.2U
M23     U115_drain ENN     U115_source VDD     P   L=.185U      W=1.4U
+  PS=.750U PD=.750U
M24     U115_source D       DmN     VDD     P   L=.185U      W=1.4U
+  PS=.750U PD=.750U
M25     VDD     U108_gate U115_drain VDD     P   L=.185U      W=1.4U
+  PS=.750U
M26     VDD     U108_gate U117_source VDD     P   L=.185U      W=1.4U
+  PS=.750U
M27     U117_source U118_gate U118_source VDD     P   L=.185U   W=1.4U
+    PS=.750U PD=.750U
M28     U118_source U122_gate DmN     VDD     P   L=.18U      W=1.57U
+  PS=.750U PD=.750U
M29     VDD     U120_gate U109_source VDD     P   L=.18U      W=1.44U
+  PS=.750U
M30     U109_source SD      DmN     VDD     P   L=.18U       W=1.44U
+  PS=.750U PD=.750U
M31     U121_drain ENN     U121_source VSS     N   L=.18U      W=0.72U
+  PS=.500U PD=.500U
M32     DmN     U122_gate U121_drain VSS     N   L=.18U      W=0.83U
+  PS=.500U PD=.500U
M33     U121_source U120_gate VSS     VSS     N   L=.18U      W=0.69U
+  PD=.500U
M34     DmN     D       U106_source VSS     N   L=.18U      W=0.69U
+  PS=.500U PD=.500U
M35     U104_drain U120_gate VSS     VSS     N   L=.18U      W=0.69U
+  PD=.500U
M36     U106_source U118_gate U104_drain VSS     N   L=.18U     W=0.69U
+   PS=.500U PD=.500U
M37     U103_drain U108_gate VSS     VSS     N   L=.18U      W=0.71U
+  PD=.500U
M38     DmN     SD      U103_drain VSS     N   L=.18U      W=0.71U
+  PS=.500U PD=.500U
M39     DmN     U15_GB  QmN     VDD     P   L=.18U      W=1.08U
+  PD=.750U
M40     DmN     U125_out QmN     VSS     N   L=.18U      W=1.04U
+  PD=.500U
M41     U128_out U125_out QmN     VDD     P   L=.187U     W=1.08U
M42     U128_out U15_GB  QmN     VSS     N   L=.18U      W=0.83U
M43     U128_in U125_out Qsl     VDD     P   L=.18U     W=1.08U
M44     U128_in U15_GB  Qsl     VSS     N   L=.18U     W=0.69U
M45     U122_gate U15_GB  Qsl     VDD     P   L=.18U     W=1.08U
M46     U122_gate U125_out Qsl     VSS     N   L=.18U    W=0.69U

.ENDS senrb4

.SUBCKT senrq4 Q  CP D ENN SC SD VDD VSS
M1      U128_out U128_in VSS     VSS     N   L=0.18U      W=0.83U
M2      U128_out U128_in VDD     VDD     P   L=0.184U      W=1.73U
M3      U128_in QmN     VSS     VSS     N   L=0.18U      W=0.83U
M4      U128_in QmN     VDD     VDD     P   L=0.184U      W=1.73U
M5      U125_out CP      VSS     VSS     N   L=0.18U      W=0.69U
M6      U125_out CP      VDD     VDD     P   L=0.184U      W=1.77U
M7      U118_gate ENN     VSS     VSS     N   L=0.18U      W=0.72U
M8      U118_gate ENN     VDD     VDD     P   L=0.18U      W=1.68U
M9      U120_gate SC      VSS     VSS     N   L=0.18U      W=0.69U
M10     U120_gate SC      VDD     VDD     P   L=0.184U      W=1.76U
M11     U108_gate U120_gate VSS     VSS     N   L=0.18U      W=0.69U
M12     U108_gate U120_gate VDD     VDD     P   L=0.18U      W=1.76U
M13     U15_GB  U125_out VSS     VSS     N   L=0.18U      W=0.68U
M14     U15_GB  U125_out VDD     VDD     P   L=0.18U      W=1.25U
M15     U122_gate U23_in  VSS     VSS     N   L=0.18U      W=0.83U
M16     U122_gate U23_in  VDD     VDD     P   L=0.184U      W=2.22U
M17     U23_in  Qsl     VSS     VSS     N   L=0.18U      W=0.83U
M18     U23_in  Qsl     VDD     VDD     P   L=0.184U      W=2.22U
M19     Q       U23_in  VSS     VSS     N   L=0.182333U      W=2.94U
M20     Q       U23_in  VDD     VDD     P   L=0.182U      W=8.2U
M21     U115_drain ENN     U115_source VDD     P   L=0.185U       W=1.40U
+  PS=.750U PD=.750U
M22     U115_source D       DmN     VDD     P   L=0.185U       W=1.40U
+  PS=.750U PD=.750U
M23     VDD     U108_gate U115_drain VDD     P   L=0.185U       W=1.40U
+  PS=.750U
M24     VDD     U108_gate U117_source VDD     P   L=0.185U       W=1.40U
+  PS=.750U
M25     U117_source U118_gate U118_source VDD     P   L=0.185U     W=1.40U
+    PS=.750U PD=.750U
M26     U118_source U122_gate DmN     VDD     P   L=0.18U       W=1.57U
+  PS=.750U PD=.750U
M27     VDD     U120_gate U109_source VDD     P   L=0.18U       W=1.44U
+  PS=.750U
M28     U109_source SD      DmN     VDD     P   L=0.18U       W=1.44U
+  PS=.750U PD=.750U
M29     U121_drain ENN     U121_source VSS     N   L=0.18U       W=0.72U
+  PS=.500U PD=.500U
M30     DmN     U122_gate U121_drain VSS     N   L=0.18U       W=0.83U
+  PS=.500U PD=.500U
M31     U121_source U120_gate VSS     VSS     N   L=0.18U       W=0.69U
+  PD=.500U
M32     DmN     D       U106_source VSS     N   L=0.18U       W=0.69U
+  PS=.500U PD=.500U
M33     U104_drain U120_gate VSS     VSS     N   L=0.18U       W=0.69U
+  PD=.500U
M34     U106_source U118_gate U104_drain VSS     N   L=0.18U      W=0.69U
+   PS=.500U PD=.500U
M35     U103_drain U108_gate VSS     VSS     N   L=0.18U       W=0.71U
+  PD=.500U
M36     DmN     SD      U103_drain VSS     N   L=0.18U       W=0.71U
+  PS=.500U PD=.500U
M37     DmN     U15_GB  QmN     VDD     P   L=0.187U       W=1.08U
+  PD=.750U
M38     DmN     U125_out QmN     VSS     N   L=0.18U       W=1.04U
+  PD=.500U
M39     U128_out U125_out QmN     VDD     P   L=0.187U      W=1.08U
M40     U128_out U15_GB  QmN     VSS     N   L=0.18U      W=0.83U
M41     U128_in U125_out Qsl     VDD     P   L=0.18U      W=1.08U
M42     U128_in U15_GB  Qsl     VSS     N   L=0.18U      W=0.69U
M43     U122_gate U15_GB  Qsl     VDD     P   L=0.18U      W=1.08U
M44     U122_gate U125_out Qsl     VSS     N   L=0.18U      W=0.69U

.ENDS senrq4

.SUBCKT sepfq1 Q  CPN D ENN SC SD SDN VDD VSS
M1      u7_S    u7_GB   QmN     VDD     P   L=0.186U         W=1.36U
M2      u7_S    u7_G    QmN     VSS     N   L=0.18U         W=0.82U
M3      DmN     u7_G    QmN     VDD     P   L=0.18U         W=1.36U
+  PD=.750U
M4      DmN     u7_GB   QmN     VSS     N   L=0.18U         W=0.68U
+  PD=.500U
M5      U130_out u7_GB   U22_in  VDD     P   L=0.187U        W=1.08U
M6      U130_out u7_G    U22_in  VSS     N   L=0.18U        W=0.55U
M7      U122_gate u7_G    U22_in  VDD     P   L=0.187U       W=1.08U
M8      U122_gate u7_GB   U22_in  VSS     N   L=0.18U       W=0.55U
M9      u7_GB   u7_G    VSS     VSS     N   L=0.18U         W=0.84U
M10     u7_GB   u7_G    VDD     VDD     P   L=0.184U         W=1.92U
M11     u7_G    CPN     VSS     VSS     N   L=0.18U         W=0.83U
M12     u7_G    CPN     VDD     VDD     P   L=0.184U         W=1.99U
M13     U116_gate ENN     VSS     VSS     N   L=0.18U       W=0.72U
M14     U116_gate ENN     VDD     VDD     P   L=0.185U       W=1.68U
M15     U120_gate SC      VSS     VSS     N   L=0.18U       W=0.83U
M16     U120_gate SC      VDD     VDD     P   L=0.184U       W=2.08U
M17     U117_gate U120_gate VSS     VSS     N   L=0.18U     W=0.71U
M18     U117_gate U120_gate VDD     VDD     P   L=0.184U     W=2.08U
M19     U22_out U22_in  VSS     VSS     N   L=0.18U         W=0.62U
M20     U22_out U22_in  VDD     VDD     P   L=0.185U         W=1.56U
M21     Q       U22_out VSS     VSS     N   L=0.18U         W=0.69U
M22     Q       U22_out VDD     VDD     P   L=0.184U         W=2.05U
M23     u7_S    U130_out VSS     VSS     N   L=0.18U        W=0.82U
M24     u7_S    U130_out VDD     VDD     P   L=0.183U        W=1.66U
M25     U116_drain U116_gate U116_source VSS     N   L=0.18U       W=0.69U
+   PS=.500U PD=.500U
M26     U121_drain ENN     U121_source VSS     N   L=0.18U         W=0.76U
+  PS=.500U PD=.500U
M27     DmN     U122_gate U121_drain VSS     N   L=0.18U           W=0.83U
+  PS=.500U PD=.500U
M28     U121_source U120_gate VSS     VSS     N   L=0.18U          W=0.83U
+  PD=.500U
M29     U116_source U120_gate VSS     VSS     N   L=0.18U          W=0.69U
+  PD=.500U
M30     DmN     D       U116_drain VSS     N   L=0.18U             W=0.69U
+  PS=.500U PD=.500U
M31     DmN     SD      U105_source VSS     N   L=0.18U            W=0.71U
+  PS=.500U PD=.500U
M32     U105_source U117_gate VSS     VSS     N   L=0.18U          W=0.71U
+  PD=.500U
M33     VDD     U117_gate U117_source VDD     P   L=0.185U          W=1.45U
+  PS=.750U
M34     U119_drain U122_gate DmN     VDD     P   L=0.185U           W=1.45U
+  PS=.750U PD=.750U
M35     U117_source U116_gate U119_drain VDD     P   L=0.185U       W=1.45U
+   PS=.750U PD=.750U
M36     VDD     U120_gate U109_source VDD     P   L=0.18U          W=1.44U
+  PS=.750U
M37     U109_source SD      DmN     VDD     P   L=0.186U            W=1.30U
+  PS=.750U PD=.750U
M38     U107_drain D       DmN     VDD     P   L=0.184U             W=1.74U
+  PS=.750U PD=.750U
M39     U115_drain ENN     U107_drain VDD     P   L=0.184U          W=1.74U
+  PS=.750U PD=.750U
M40     VDD     U117_gate U115_drain VDD     P   L=0.18U           W=1.40U
+  PS=.750U
M41     U130_out SDN     VDD     VDD     P   L=0.185U               W=1.53U
M42     U130_out QmN     VDD     VDD     P   L=0.187U               W=1.14U
M43     U130_$$7 SDN     VSS     VSS     N   L=0.18U               W=0.75U
M44     U130_out QmN     U130_$$7 VSS     N   L=0.18U              W=0.75U
M45     U122_gate SDN     VDD     VDD     P   L=0.185U              W=1.45U
M46     U122_gate U22_out VDD     VDD     P   L=0.185U              W=1.45U
M47     U129_$$7 SDN     VSS     VSS     N   L=0.18U               W=0.83U
M48     U122_gate U22_out U129_$$7 VSS     N   L=0.18U             W=0.83U

.ENDS sepfq1

.SUBCKT sepfq2 Q  CPN D ENN SC SD SDN VDD VSS
M1      u7_S    u7_GB   QmN     VDD     P   L=.186U  W=1.36U  
M2      u7_S    u7_G    QmN     VSS     N   L=.180U  W=0.82U  
M3      DmN     u7_G    QmN     VDD     P   L=.180U  W=1.36U   
+  PD=.750U
M4      DmN     u7_GB   QmN     VSS     N   L=.180U  W=0.68U   PD=.500U
M5      U130_out u7_GB   U22_in  VDD     P   L=.187U  W=1.08U  
M6      U130_out u7_G    U22_in  VSS     N   L=.180U  W=0.55U  
M7      U122_gate u7_G    U22_in  VDD     P   L=.180U  W=1.08U  
M8      U122_gate u7_GB   U22_in  VSS     N   L=.180U  W=0.55U  
M9      u7_GB   u7_G    VSS     VSS     N   L=.180U  W=0.84U  
M10     u7_GB   u7_G    VDD     VDD     P   L=.180U  W=1.92U  
M11     u7_G    CPN     VSS     VSS     N   L=.180U  W=0.83U  
M12     u7_G    CPN     VDD     VDD     P   L=.184U  W=1.99U  
M13     U116_gate ENN     VSS     VSS     N   L=.180U  W=0.72U  
M14     U116_gate ENN     VDD     VDD     P   L=.180U  W=1.68U  
M15     U120_gate SC      VSS     VSS     N   L=.180U  W=0.83U  
M16     U120_gate SC      VDD     VDD     P   L=.184U  W=2.08U  
M17     U117_gate U120_gate VSS     VSS     N   L=.180U  W=0.71U  
M18     U117_gate U120_gate VDD     VDD     P   L=.180U  W=2.08U  
M19     U22_out U22_in  VSS     VSS     N   L=.180U  W=0.62U  
M20     U22_out U22_in  VDD     VDD     P   L=.180U  W=1.5U  
M21     Q       U22_out VSS     VSS     N   L=.185U  W=1.43U  
M22     Q       U22_out VDD     VDD     P   L=.184U  W=4.1U  
M23     u7_S    U130_out VSS     VSS     N   L=.180U  W=0.82U  
M24     u7_S    U130_out VDD     VDD     P   L=.185U  W=1.66U  
M25     U116_drain U116_gate U116_source VSS     N   L=.180U  W=0.69U  
+   PS=.500U PD=.500U
M26     U121_drain ENN     U121_source VSS     N   L=.180U  W=0.76U   
+  PS=.500U PD=.500U
M27     DmN     U122_gate U121_drain VSS     N   L=.180U  W=0.83U   
+  PS=.500U PD=.500U
M28     U121_source U120_gate VSS     VSS     N   L=.180U  W=0.83U   
+  PD=.500U
M29     U116_source U120_gate VSS     VSS     N   L=.180U  W=0.69U   
+  PD=.500U
M30     DmN     D       U116_drain VSS     N   L=.180U  W=0.69U   
+  PS=.500U PD=.500U
M31     DmN     SD      U105_source VSS     N   L=.180U  W=0.71U   
+  PS=.500U PD=.500U
M32     U105_source U117_gate VSS     VSS     N   L=.180U  W=0.71U   
+  PD=.500U
M33     VDD     U117_gate U117_source VDD     P   L=.180U  W=1.45U   
+  PS=.750U
M34     U119_drain U122_gate DmN     VDD     P   L=.185U  W=1.45U   
+  PS=.750U PD=.750U
M35     U117_source U116_gate U119_drain VDD     P   L=.185U  W=1.45U  
+   PS=.750U PD=.750U
M36     VDD     U120_gate U109_source VDD     P   L=.186U  W=1.44U   
+  PS=.750U
M37     U109_source SD      DmN     VDD     P   L=.186U  W=1.3U   
+  PS=.750U PD=.750U
M38     U107_drain D       DmN     VDD     P   L=.180U  W=1.74U   
+  PS=.750U PD=.750U
M39     U115_drain ENN     U107_drain VDD     P   L=.180U  W=1.74U   
+  PS=.750U PD=.750U
M40     VDD     U117_gate U115_drain VDD     P   L=.185U  W=1.4U   
+  PS=.750U
M41     U130_out SDN     VDD     VDD     P   L=.185U  W=1.53U  
M42     U130_out QmN     VDD     VDD     P   L=.180U  W=1.14U  
M43     U130_$$7 SDN     VSS     VSS     N   L=.180U  W=0.75U  
M44     U130_out QmN     U130_$$7 VSS     N   L=.180U  W=0.75U  
M45     U122_gate SDN     VDD     VDD     P   L=.185U  W=1.45U  
M46     U122_gate U22_out VDD     VDD     P   L=.186U  W=1.45U  
M47     U129_$$7 SDN     VSS     VSS     N   L=.180U  W=0.83U  
M48     U122_gate U22_out U129_$$7 VSS     N   L=.180U  W=0.83U  

.ENDS sepfq2

.SUBCKT sepfq4 Q  CPN D ENN SC SD SDN VDD VSS
M1      u7_S    u7_GB   QmN     VDD     P   L=0.186U  W=1.36U  
M2      u7_S    u7_G    QmN     VSS     N   L=0.180U  W=0.82U  
M3      DmN     u7_G    QmN     VDD     P   L=0.180U  W=1.36U   
+  PD=.750U
M4      DmN     u7_GB   QmN     VSS     N   L=0.180U  W=0.68U   PD=.500U
M5      U130_out u7_GB   U22_in  VDD     P   L=0.187U  W=1.08U  
M6      U130_out u7_G    U22_in  VSS     N   L=0.180U  W=0.55U  
M7      U122_gate u7_G    U22_in  VDD     P   L=0.180U  W=1.08U  
M8      U122_gate u7_GB   U22_in  VSS     N   L=0.180U  W=0.55U  
M9      u7_GB   u7_G    VSS     VSS     N   L=0.180U  W=0.84U  
M10     u7_GB   u7_G    VDD     VDD     P   L=0.180U  W=1.92U  
M11     u7_G    CPN     VSS     VSS     N   L=0.180U  W=0.83U  
M12     u7_G    CPN     VDD     VDD     P   L=0.184U  W=1.99U  
M13     U116_gate ENN     VSS     VSS     N   L=0.180U  W=0.72U  
M14     U116_gate ENN     VDD     VDD     P   L=0.180U  W=1.68U  
M15     U120_gate SC      VSS     VSS     N   L=0.180U  W=0.83U  
M16     U120_gate SC      VDD     VDD     P   L=0.185U  W=2.08U  
M17     U117_gate U120_gate VSS     VSS     N   L=0.180U  W=0.71U  
M18     U117_gate U120_gate VDD     VDD     P   L=0.180U  W=2.08U  
M19     U22_out U22_in  VSS     VSS     N   L=0.180U  W=0.93U  
M20     U22_out U22_in  VDD     VDD     P   L=0.180U  W=2.05U  
M21     Q       U22_out VSS     VSS     N   L=0.180U  W=2.78U  
M22     Q       U22_out VDD     VDD     P   L=0.183U  W=8.2U  
M23     u7_S    U130_out VSS     VSS     N   L=0.180U  W=0.82U  
M24     u7_S    U130_out VDD     VDD     P   L=0.185U  W=1.66U  
M25     U116_drain U116_gate U116_source VSS     N   L=0.180U  W=0.69U  
+   PS=.500U PD=.500U
M26     U121_drain ENN     U121_source VSS     N   L=0.180U  W=0.76U   
+  PS=.500U PD=.500U
M27     DmN     U122_gate U121_drain VSS     N   L=0.180U  W=0.83U   
+  PS=.500U PD=.500U
M28     U121_source U120_gate VSS     VSS     N   L=0.180U  W=0.83U   
+  PD=.500U
M29     U116_source U120_gate VSS     VSS     N   L=0.180U  W=0.69U   
+  PD=.500U
M30     DmN     D       U116_drain VSS     N   L=0.180U  W=0.69U   
+  PS=.500U PD=.500U
M31     DmN     SD      U105_source VSS     N   L=0.180U  W=0.71U   
+  PS=.500U PD=.500U
M32     U105_source U117_gate VSS     VSS     N   L=0.180U  W=0.71U   
+  PD=.500U
M33     VDD     U117_gate U117_source VDD     P   L=0.180U  W=1.45U   
+  PS=.750U
M34     U119_drain U122_gate DmN     VDD     P   L=0.185U  W=1.45U   
+  PS=.750U PD=.750U
M35     U117_source U116_gate U119_drain VDD     P   L=0.185U  W=1.45U  
+   PS=.750U PD=.750U
M36     VDD     U120_gate U109_source VDD     P   L=0.186U  W=1.44U   
+  PS=.750U
M37     U109_source SD      DmN     VDD     P   L=0.186U  W=1.3U   
+  PS=.750U PD=.750U
M38     U107_drain D       DmN     VDD     P   L=0.180U  W=1.74U   
+  PS=.750U PD=.750U
M39     U115_drain ENN     U107_drain VDD     P   L=0.180U  W=1.74U   
+  PS=.750U PD=.750U
M40     VDD     U117_gate U115_drain VDD     P   L=0.185U  W=1.4U   
+  PS=.750U
M41     U130_out SDN     VDD     VDD     P   L=0.185U  W=1.53U  
M42     U130_out QmN     VDD     VDD     P   L=0.180U  W=1.14U  
M43     U130_$$7 SDN     VSS     VSS     N   L=0.180U  W=0.75U  
M44     U130_out QmN     U130_$$7 VSS     N   L=0.180U  W=0.75U  
M45     U122_gate SDN     VDD     VDD     P   L=0.185U  W=1.45U  
M46     U122_gate U22_out VDD     VDD     P   L=0.185U  W=1.45U  
M47     U129_$$7 SDN     VSS     VSS     N   L=0.180U  W=0.83U  
M48     U122_gate U22_out U129_$$7 VSS     N   L=0.180U  W=0.83U  

.ENDS sepfq4

.SUBCKT seprq4 Q  CP D ENN SC SD SDN VDD VSS
M1      DmN     U15_GB  QmN     VDD     P   L=0.186U  W=1.36U   
+  PD=.750U
M2      DmN     U15_G   QmN     VSS     N   L=0.18U  W=0.68U   PD=.500U
M3      u7_S    U15_G   QmN     VDD     P   L=0.18U  W=1.36U  
M4      u7_S    U15_GB  QmN     VSS     N   L=0.18U  W=0.82U  
M5      U130_out U15_G   U22_in  VDD     P   L=0.18U  W=1.08U  
M6      U130_out U15_GB  U22_in  VSS     N   L=0.18U  W=0.55U  
M7      U119_gate U15_GB  U22_in  VDD     P   L=0.18U  W=1.08U  
M8      U119_gate U15_G   U22_in  VSS     N   L=0.18U  W=0.55U  
M9      U15_GB  U15_G   VSS     VSS     N   L=0.18U  W=0.84U  
M10     U15_GB  U15_G   VDD     VDD     P   L=0.18U  W=1.92U  
M11     U15_G   CP      VSS     VSS     N   L=0.18U  W=0.83U  
M12     U15_G   CP      VDD     VDD     P   L=0.184U  W=1.99U  
M13     U118_gate ENN     VSS     VSS     N   L=0.18U  W=0.72U  
M14     U118_gate ENN     VDD     VDD     P   L=0.185U  W=1.68U  
M15     U120_gate SC      VSS     VSS     N   L=0.18U  W=0.83U  
M16     U120_gate SC      VDD     VDD     P   L=0.184U  W=2.08U  
M17     U117_gate U120_gate VSS     VSS     N   L=0.18U  W=0.71U  
M18     U117_gate U120_gate VDD     VDD     P   L=0.184U  W=2.08U  
M19     U22_out U22_in  VSS     VSS     N   L=0.18U  W=0.93U  
M20     U22_out U22_in  VDD     VDD     P   L=0.184U  W=2.05U  
M21     Q       U22_out VSS     VSS     N   L=0.18U  W=2.78U  
M22     Q       U22_out VDD     VDD     P   L=0.183U  W=8.2U  
M23     u7_S    U130_out VSS     VSS     N   L=0.18U  W=0.82U  
M24     u7_S    U130_out VDD     VDD     P   L=0.185U  W=1.59U  
M25     U119_drain U119_gate DmN     VDD     P   L=0.18U  W=1.45U   
+  PS=.750U PD=.750U
M26     U118_drain U118_gate U119_drain VDD     P   L=0.18U  W=1.45U   
+  PS=.750U PD=.750U
M27     VDD     U117_gate U118_drain VDD     P   L=0.18U  W=1.45U   
+  PS=.750U
M28     VDD     U120_gate U109_source VDD     P   L=0.18U  W=1.44U   
+  PS=.750U
M29     U109_source SD      DmN     VDD     P   L=0.186U  W=1.3U   
+  PS=.750U PD=.750U
M30     U107_drain D       DmN     VDD     P   L=0.185U  W=1.74U   
+  PS=.750U PD=.750U
M31     U115_drain ENN     U107_drain VDD     P   L=0.185U  W=1.74U   
+  PS=.750U PD=.750U
M32     VDD     U117_gate U115_drain VDD     P   L=0.18U  W=1.4U   
+  PS=.750U
M33     U120_drain U120_gate VSS     VSS     N   L=0.18U  W=0.83U   
+  PD=.500U
M34     U104_drain U120_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.500U
M35     DmN     D       U106_source VSS     N   L=0.18U  W=0.69U   
+  PS=.500U PD=.500U
M36     DmN     U119_gate U122_source VSS     N   L=0.18U  W=0.83U   
+  PS=.500U PD=.500U
M37     U122_source ENN     U120_drain VSS     N   L=0.18U  W=0.76U   
+  PS=.500U PD=.500U
M38     U106_source U118_gate U104_drain VSS     N   L=0.18U  W=0.69U  
+   PS=.500U PD=.500U
M39     DmN     SD      U105_source VSS     N   L=0.18U  W=0.71U   
+  PS=.500U PD=.500U
M40     U105_source U117_gate VSS     VSS     N   L=0.18U  W=0.71U   
+  PD=.500U
M41     U130_out SDN     VDD     VDD     P   L=0.18U  W=1.52U  
M42     U130_out QmN     VDD     VDD     P   L=0.188U  W=1.13U  
M43     U130_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.75U  
M44     U130_out QmN     U130_$$7 VSS     N   L=0.18U  W=0.75U  
M45     U119_gate SDN     VDD     VDD     P   L=0.186U  W=1.45U  
M46     U119_gate U22_out VDD     VDD     P   L=0.18U  W=1.45U  
M47     U129_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.83U 
M48     U119_gate U22_out U129_$$7 VSS     N   L=0.18U  W=0.83U  

.ENDS seprq4

.SUBCKT skbrb1 Q QN  CP CDN J KZ SC SD SDN VDD VSS
M1      u7_S    u7_GB   u7_D    VDD     P   L=0.18U  PD=.750U  W=1.29U
M2      u7_S    u7_G    u7_D    VSS     N   L=0.18U  PD=.750U  W=0.55U
M3      U15_S   u7_G    u7_D    VDD     P   L=0.186U  PD=.797U  W=1.43U
M4      U15_S   u7_GB   u7_D    VSS     N   L=0.18U  PD=.600U  W=0.50U
M5      U24_out u7_GB   u8_D    VDD     P   L=0.18U  PD=.900U  W=1.08U
M6      U24_out u7_G    u8_D    VSS     N   L=0.18U  W=0.42U
+  PD=1.045U
M7      U77_gate u7_G    u8_D    VDD     P   L=0.18U  W=0.75U
+  PD=.705U
M8      U77_gate u7_GB   u8_D    VSS     N   L=0.18U  W=0.42U
+  PD=.920U
M9      u7_G    u7_GB   VSS     VSS     N   L=0.18U  W=0.35U
M10     u7_G    u7_GB   VDD     VDD     P   L=0.18U  W=1.08U
M11     Q       U21_in  VSS     VSS     N   L=0.18U  W=0.69U
M12     Q       U21_in  VDD     VDD     P   L=0.184U  W=2.05U
M13     u7_GB   CP      VSS     VSS     N   L=0.18U  W=0.35U
M14     u7_GB   CP      VDD     VDD     P   L=0.18U  W=1.0U
M15     U75_gate U77_gate VSS     VSS     N   L=0.18U  W=0.58U
M16     U75_gate U77_gate VDD     VDD     P   L=0.18U  W=1.49U
M17     U90_gate SC      VSS     VSS     N   L=0.18U  W=0.26U
M18     U90_gate SC      VDD     VDD     P   L=0.18U  W=0.88U
M19     U92_gate U90_gate VSS     VSS     N   L=0.18U  W=0.36U
M20     U92_gate U90_gate VDD     VDD     P   L=0.18U  W=1.30U
M21     QN      u8_D    VSS     VSS     N   L=0.18U  W=0.69U
M22     QN      u8_D    VDD     VDD     P   L=0.184U  W=2.05U
M23     U15_S   U92_gate U92_source VSS     N   L=0.18U  W=0.76U
+  PS=.300U PD=.600U
M24     U76_drain KZ      U15_S   VSS     N   L=0.18U  W=1.04U
+  PS=.600U PD=.750U
M25     U90_drain U90_gate VSS     VSS     N   L=0.18U  W=0.36U
+  PD=.600U
M26     U76_drain U77_gate U90_drain VSS     N   L=0.18U  W=1.04U
+  PS=.600U PD=.750U
M27     U76_drain J       U90_drain VSS     N   L=0.18U  W=0.58U
+  PS=.600U PD=.750U
M28     U15_S   U75_gate U76_drain VSS     N   L=0.18U  W=0.58U
+  PS=.750U PD=.600U
M29     U92_source SD      VSS     VSS     N   L=0.18U  W=0.76U
+  PD=.300U
M30     U24_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.53U
+  PD=1.045U
M31     U24_out u7_D    U24_u7_drain VSS     N   L=0.18U  W=0.53U
+  PS=1.045U PD=1.045U
M32     U24_out u7_D    VDD     VDD     P   L=0.18U  PD=.900U  W=0.91U
M33     VDD     SDN     U24_out VDD     P   L=0.187U  PS=.900U  W=1.18U
M34     U81_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.73U
+  PD=1.370U
M35     U21_in  u8_D    U81_u7_drain VSS     N   L=0.18U  W=0.73U
+  PS=1.370U PD=1.370U
M36     U21_in  u8_D    VDD     VDD     P   L=0.18U  W=0.99U
+  PD=1.005U
M37     VDD     CDN     U21_in  VDD     P   L=0.187U  W=1.15U
+  PS=1.005U
M38     U82_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.73U
+  PD=.920U
M39     U77_gate U21_in  U82_u7_drain VSS     N   L=0.18U  W=0.73U
+  PS=.920U PD=.920U
M40     U77_gate U21_in  VDD     VDD     P   L=0.18U  W=0.82U
+  PD=.705U
M41     VDD     SDN     U77_gate VDD     P   L=0.18U  W=0.82U
+  PS=.705U
M42     U80_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.73U
+  PD=.750U
M43     u7_S    U24_out U80_u7_drain VSS     N   L=0.18U  W=0.73U
+  PS=.750U PD=.750U
M44     u7_S    U24_out VDD     VDD     P   L=0.187U  PD=.750U  W=1.18U
M45     VDD     CDN     u7_S    VDD     P   L=0.187U  PS=.750U  W=1.18U
M46     U15_S   KZ      U73_source VDD     P   L=0.18U  W=1.47U
+  PS=1.045U PD=.797U
M47     U73_source U75_gate U72_source VDD     P   L=0.18U  W=1.47U
+  PS=.797U PD=1.045U
M48     U72_source U77_gate U74_source VDD     P   L=0.18U  W=1.47U
+  PS=1.045U PD=.797U
M49     U74_source J       U15_S   VDD     P   L=0.18U  W=1.47U
+  PS=.797U PD=1.045U
M50     U72_source U92_gate VDD     VDD     P   L=0.186U  W=1.38U
+  PD=.797U
M51     U15_S   U90_gate U94_source VDD     P   L=0.18U  W=1.52U
+  PS=.300U PD=.797U
M52     U94_source SD      VDD     VDD     P   L=0.18U  W=1.52U
+  PD=.300U

.ENDS skbrb1

.SUBCKT skbrb2 Q QN  CP CDN J KZ SC SD SDN VDD VSS
M1      u7_S    u7_GB   u7_D    VDD     P   L=0.18U  PD=.750U  W=1.29U
M2      u7_S    u7_G    u7_D    VSS     N   L=0.18U  PD=.750U  W=0.55U
M3      U15_S   u7_G    u7_D    VDD     P   L=0.186U  PD=.797U  W=1.43U
M4      U15_S   u7_GB   u7_D    VSS     N   L=0.18U  PD=.600U  W=0.5U
M5      u8_S    u7_GB   U81_in1 VDD     P   L=0.18U  PD=.900U  W=1.08U
M6      u8_S    u7_G    U81_in1 VSS     N   L=0.18U  W=0.42U
+  PD=1.045U
M7      U77_gate u7_G    U81_in1 VDD     P   L=0.18U  W=0.75U
+  PD=.705U
M8      U77_gate u7_GB   U81_in1 VSS     N   L=0.18U  W=0.42U
+  PD=.920U
M9      u7_G    u7_GB   VSS     VSS     N   L=0.18U  W=0.35U
M10     u7_G    u7_GB   VDD     VDD     P   L=0.18U  W=1.08U
M11     Q       U81_out VSS     VSS     N   L=0.18U  W=1.45U
M12     Q       U81_out VDD     VDD     P   L=0.184U W=4.1U
M13     u7_GB   CP      VSS     VSS     N   L=0.18U  W=0.35U
M14     u7_GB   CP      VDD     VDD     P   L=0.18U  W=1.0U
M15     U75_gate U77_gate VSS     VSS     N   L=0.18U  W=0.58U
M16     U75_gate U77_gate VDD     VDD     P   L=0.18U W=1.49U
M17     U90_gate SC      VSS     VSS     N   L=0.18U  W=0.26U
M18     U90_gate SC      VDD     VDD     P   L=0.18U  W=0.88U
M19     U92_gate U90_gate VSS     VSS     N   L=0.18U  W=0.36U
M20     U92_gate U90_gate VDD     VDD     P   L=0.18U  W=1.3U
M21     QN      U81_in1 VSS     VSS     N   L=0.18U  W=1.45U
M22     QN      U81_in1 VDD     VDD     P   L=0.184U W=4.1U
M23     U81_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.73U
+  PD=1.370U
M24     U81_out U81_in1 U81_u7_drain VSS     N   L=0.18U  W=0.73U
+  PS=1.370U PD=1.370U
M25     U81_out U81_in1 VDD     VDD     P   L=0.18U  W=0.99U
+  PD=1.005U
M26     VDD     CDN     U81_out VDD     P   L=0.187U  W=1.15U
+  PS=1.005U
M27     U24_u7_drain SDN     VSS     VSS     N   L=0.18U W=0.53U
+  PD=1.045U
M28     u8_S    u7_D    U24_u7_drain VSS     N   L=0.18U W=0.53U
+  PS=1.045U PD=1.045U
M29     u8_S    u7_D    VDD     VDD     P   L=0.18U  PD=.900U  W=0.91U
M30     VDD     SDN     u8_S    VDD     P   L=0.187U  PS=.900U  W=1.18U
M31     U82_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.73U
+  PD=.920U
M32     U77_gate U81_out U82_u7_drain VSS     N   L=0.18U  W=0.73U
+  PS=.920U PD=.920U
M33     U77_gate U81_out VDD     VDD     P   L=0.18U  W=0.82U
+  PD=.705U
M34     VDD     SDN     U77_gate VDD     P   L=0.18U  W=0.82U
+  PS=.705U
M35     U80_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.73U
+  PD=.750U
M36     u7_S    u8_S    U80_u7_drain VSS     N   L=0.18U  W=0.73U
+  PS=.750U PD=.750U
M37     u7_S    u8_S    VDD     VDD     P   L=0.187U  PD=.750U  W=1.18U
M38     VDD     CDN     u7_S    VDD     P   L=0.187U  PS=.750U  W=1.18U
M39     U15_S   U92_gate U92_source VSS     N   L=0.18U  W=0.76U
+  PS=.300U PD=.600U
M40     U76_drain KZ      U15_S   VSS     N   L=0.18U  W=1.04U
+  PS=.600U PD=.750U
M41     U90_drain U90_gate VSS     VSS     N   L=0.18U  W=0.36U
+  PD=.600U
M42     U76_drain U77_gate U90_drain VSS     N   L=0.18U  W=1.04U
+  PS=.600U PD=.750U
M43     U76_drain J       U90_drain VSS     N   L=0.18U  W=0.58U
+  PS=.600U PD=.750U
M44     U15_S   U75_gate U76_drain VSS     N   L=0.18U  W=0.58U
+  PS=.750U PD=.600U
M45     U92_source SD      VSS     VSS     N   L=0.18U  W=0.76U
+  PD=.300U
M46     U15_S   KZ      U73_source VDD     P   L=0.18U  W=1.47U
+  PS=1.045U PD=.797U
M47     U73_source U75_gate U72_source VDD     P   L=0.18U  W=1.47U
+  PS=.797U PD=1.045U
M48     U72_source U77_gate U74_source VDD     P   L=0.18U  W=1.47U
+  PS=1.045U PD=.797U
M49     U74_source J       U15_S   VDD     P   L=0.18U  W=1.47U
+  PS=.797U PD=1.045U
M50     U72_source U92_gate VDD     VDD     P   L=0.186U  W=1.38U
+  PD=.797U
M51     U15_S   U90_gate U94_source VDD     P   L=0.18U  W=1.52U
+  PS=.300U PD=.797U
M52     U94_source SD      VDD     VDD     P   L=0.18U  W=1.52U
+  PD=.300U

.ENDS skbrb2

.SUBCKT skbrb4 Q QN  CP CDN J KZ SC SD SDN VDD VSS
M1      u7_S    u7_GB   u7_D    VDD     P   L=0.18U  PD=.750U  W=1.29U
M2      u7_S    u7_G    u7_D    VSS     N   L=0.18U  PD=.750U  W=0.55U
M3      U15_S   u7_G    u7_D    VDD     P   L=0.186U  PD=.797U  W=1.43U
M4      U15_S   u7_GB   u7_D    VSS     N   L=0.18U  PD=.600U  W=0.5U
M5      u8_S    u7_GB   U81_in1 VDD     P   L=0.18U  PD=.900U  W=1.08U
M6      u8_S    u7_G    U81_in1 VSS     N   L=0.18U  W=0.42U
+  PD=1.045U
M7      U77_gate u7_G    U81_in1 VDD     P   L=0.18U  W=0.75U
+  PD=.705U
M8      U77_gate u7_GB   U81_in1 VSS     N   L=0.18U  W=0.42U
+  PD=.920U
M9      u7_G    u7_GB   VSS     VSS     N   L=0.18U  W=0.35U
M10     u7_G    u7_GB   VDD     VDD     P   L=0.18U  W=1.08U
M11     Q       U81_out VSS     VSS     N   L=0.18U  W=2.94U
M12     Q       U81_out VDD     VDD     P   L=0.184U  W=8.2U
M13     u7_GB   CP      VSS     VSS     N   L=0.18U  W=0.35U
M14     u7_GB   CP      VDD     VDD     P   L=0.18U  W=1.0U
M15     U75_gate U77_gate VSS     VSS     N   L=0.18U  W=0.58U
M16     U75_gate U77_gate VDD     VDD     P   L=0.18U  W=1.49U
M17     U90_gate SC      VSS     VSS     N   L=0.18U  W=0.26U
M18     U90_gate SC      VDD     VDD     P   L=0.18U  W=0.88U
M19     U92_gate U90_gate VSS     VSS     N   L=0.18U  W=0.36U
M20     U92_gate U90_gate VDD     VDD     P   L=0.18U  W=1.30U
M21     QN      U81_in1 VSS     VSS     N   L=0.18U  W=3.10U
M22     QN      U81_in1 VDD     VDD     P   L=0.184U  W=8.2U
M23     U81_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.73U
+  PD=1.370U
M24     U81_out U81_in1 U81_u7_drain VSS     N   L=0.18U  W=0.73U
+  PS=1.370U PD=1.370U
M25     U81_out U81_in1 VDD     VDD     P   L=0.18U  W=0.99U
+  PD=1.005U
M26     VDD     CDN     U81_out VDD     P   L=0.187U  W=1.15U
+  PS=1.005U
M27     U24_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.53U
+  PD=1.045U
M28     u8_S    u7_D    U24_u7_drain VSS     N   L=0.18U  W=0.53U
+  PS=1.045U PD=1.045U
M29     u8_S    u7_D    VDD     VDD     P   L=0.18U  PD=.900U  W=0.91U
M30     VDD     SDN     u8_S    VDD     P   L=0.187U  PS=.900U  W=1.18U
M31     U82_u7_drain SDN     VSS     VSS     N   L=0.18U  W=0.73U
+  PD=.920U
M32     U77_gate U81_out U82_u7_drain VSS     N   L=0.18U  W=0.73U
+  PS=.920U PD=.920U
M33     U77_gate U81_out VDD     VDD     P   L=0.18U  W=0.823846153846154U
+  PD=.705U
M34     VDD     SDN     U77_gate VDD     P   L=0.18U  W=0.823846153846154U
+  PS=.705U
M35     U80_u7_drain CDN     VSS     VSS     N   L=0.18U  W=0.73U
+  PD=.750U
M36     u7_S    u8_S    U80_u7_drain VSS     N   L=0.18U  W=0.73U
+  PS=.750U PD=.750U
M37     u7_S    u8_S    VDD     VDD     P   L=0.187U  PD=.750U  W=1.18U
M38     VDD     CDN     u7_S    VDD     P   L=0.187U  PS=.750U  W=1.18U
M39     U15_S   U92_gate U92_source VSS     N   L=0.18U  W=0.76U
+  PS=.300U PD=.600U
M40     U76_drain KZ      U15_S   VSS     N   L=0.18U  W=1.04U
+  PS=.600U PD=.750U
M41     U90_drain U90_gate VSS     VSS     N   L=0.18U  W=0.36U
+  PD=.600U
M42     U76_drain U77_gate U90_drain VSS     N   L=0.18U  W=1.04U
+  PS=.600U PD=.750U
M43     U76_drain J       U90_drain VSS     N   L=0.18U  W=0.58U
+  PS=.600U PD=.750U
M44     U15_S   U75_gate U76_drain VSS     N   L=0.18U  W=0.58U
+  PS=.750U PD=.600U
M45     U92_source SD      VSS     VSS     N   L=0.18U  W=0.76U
+  PD=.300U
M46     U15_S   KZ      U73_source VDD     P   L=0.18U  W=1.47U
+  PS=1.045U PD=.797U
M47     U73_source U75_gate U72_source VDD     P   L=0.18U  W=1.47U
+  PS=.797U PD=1.045U
M48     U72_source U77_gate U74_source VDD     P   L=0.18U  W=1.47U
+  PS=1.045U PD=.797U
M49     U74_source J       U15_S   VDD     P   L=0.18U  W=1.47U
+  PS=.797U PD=1.045U
M50     U72_source U92_gate VDD     VDD     P   L=0.186U  W=1.38U
+  PD=.797U
M51     U15_S   U90_gate U94_source VDD     P   L=0.18U  W=1.52U
+  PS=.300U PD=.797U
M52     U94_source SD      VDD     VDD     P   L=0.18U  W=1.52U
+  PD=.300U

.ENDS skbrb4

.SUBCKT slbhb1 SO Q QN  CDN D E SC SD SDN VDD VSS
M1      U82_out SDN     VDD     VDD     P   L=0.184444U  W=1.83U    
M2      U82_out U82_in1 VDD     VDD     P   L=0.18U  W=1.83U    
M3      U82_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.82U    
M4      U82_out U82_in1 U82_$$7 VSS     N   L=0.18U  W=0.82U    
M5      U76_out CDN     VDD     VDD     P   L=0.185U  W=1.7U    
M6      U76_out U82_out VDD     VDD     P   L=0.185U  W=1.68U    
M7      U76_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.83U    
M8      U76_out U82_out U76_$$7 VSS     N   L=0.18U  W=0.83U    
M9      U76_out u7_GB   U82_in1 VDD     P   L=0.18U  W=1.41U    
M10     U76_out u7_G    U82_in1 VSS     N   L=0.18U  W=0.46U    
M11     U48_drain u7_G    U82_in1 VDD     P   L=0.185U  W=1.41U     
+  PD=.447U
M12     U48_drain u7_GB   U82_in1 VSS     N   L=0.18U  W=0.46U     
+  PD=.480U
M13     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.82U    
M14     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.5U    
M15     U82_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.82U    
M16     U82_out u7_G    u9_D    VSS     N   L=0.18U  W=0.54U    
M17     U48_drain D       U48_source VSS     N   L=0.18U  W=0.68U     
+  PS=.480U PD=.480U
M18     U48_source U68_gate U68_source VSS     N   L=0.18U  W=0.68U     
+  PS=.420U PD=.480U
M19     U69_drain U43_gate U68_source VSS     N   L=0.18U  W=0.68U     
+  PS=.420U PD=.480U
M20     U68_source CDN     VSS     VSS     N   L=0.18U  W=0.69U     
+  PD=.420U
M21     U48_drain SD      U69_drain VSS     N   L=0.18U  W=0.68U     
+  PS=.480U PD=.480U
M22     U66_drain SD      U48_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.447U PD=.520U
M23     VDD     U68_gate U66_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.520U
M24     U67_drain D       U48_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.447U PD=.520U
M25     VDD     U43_gate U67_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.520U
M26     VDD     CDN     U48_drain VDD     P   L=0.184U  W=1.91U     
+  PS=.447U
M27     u7_G    E       VSS     VSS     N   L=0.18U  W=0.66U    
M28     u7_G    E       VDD     VDD     P   L=0.18U  W=1.54U    
M29     u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.66U    
M30     u7_GB   u7_G    VDD     VDD     P   L=0.185U  W=1.54U    
M31     U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U    
M32     U43_gate U68_gate VDD     VDD     P   L=0.18U  W=1.8U    
M33     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U    
M34     U68_gate SC      VDD     VDD     P   L=0.184U  W=1.91U    
M35     u9_S    U78_in  VSS     VSS     N   L=0.18U  W=0.83U    
M36     u9_S    U78_in  VDD     VDD     P   L=0.184U  W=1.87U    
M37     U78_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U    
M38     U78_in  u9_D    VDD     VDD     P   L=0.184U  W=1.87U    
M39     Q       U20_in  VSS     VSS     N   L=0.18U  W=0.69U    
M40     Q       U20_in  VDD     VDD     P   L=0.184U  W=2.05U    
M41     QN      U83_in  VSS     VSS     N   L=0.18U  W=0.69U    
M42     QN      U83_in  VDD     VDD     P   L=0.184U  W=2.05U    
M43     U83_in  U76_out VSS     VSS     N   L=0.18U  W=0.69U    
M44     U83_in  U76_out VDD     VDD     P   L=0.185U  W=1.76U    
M45     U20_in  U82_out VSS     VSS     N   L=0.18U  W=0.69U    
M46     U20_in  U82_out VDD     VDD     P   L=0.184U  W=2.05U    
M47     SO      U78_in  VSS     VSS     N   L=0.18U  W=0.69U    
M48     SO      U78_in  VDD     VDD     P   L=0.184U  W=2.05U    

.ENDS slbhb1

.SUBCKT slbhb2 SO Q QN  CDN D E SC SD SDN VDD VSS
M1      U82_out SDN     VDD     VDD     P   L=0.18U  W=1.83U    
M2      U82_out U82_in1 VDD     VDD     P   L=0.184U  W=1.83U    
M3      U82_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.83U    
M4      U82_out U82_in1 U82_$$7 VSS     N   L=0.18U  W=0.83U    
M5      U76_out CDN     VDD     VDD     P   L=0.185U  W=1.7U    
M6      U76_out U82_out VDD     VDD     P   L=0.185U  W=1.68U    
M7      U76_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.83U    
M8      U76_out U82_out U76_$$7 VSS     N   L=0.18U  W=0.83U    
M9      U76_out u7_GB   U82_in1 VDD     P   L=0.18U  W=1.41U    
M10     U76_out u7_G    U82_in1 VSS     N   L=0.18U  W=0.46U    
M11     U48_drain u7_G    U82_in1 VDD     P   L=0.185U  W=1.41U     
+  PD=.447U
M12     U48_drain u7_GB   U82_in1 VSS     N   L=0.18U  W=0.46U     
+  PD=.480U
M13     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.82U    
M14     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.54U    
M15     U82_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.82U    
M16     U82_out u7_G    u9_D    VSS     N   L=0.18U  W=0.54U    
M17     U48_drain D       U48_source VSS     N   L=0.18U  W=0.68U     
+  PS=.480U PD=.480U
M18     U48_source U68_gate U68_source VSS     N   L=0.18U  W=0.68U     
+  PS=.420U PD=.480U
M19     U69_drain U43_gate U68_source VSS     N   L=0.18U  W=0.68U     
+  PS=.420U PD=.480U
M20     U68_source CDN     VSS     VSS     N   L=0.18U  W=0.69U     
+  PD=.420U
M21     U48_drain SD      U69_drain VSS     N   L=0.18U  W=0.68U     
+  PS=.480U PD=.480U
M22     U66_drain SD      U48_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.447U PD=.520U
M23     VDD     U68_gate U66_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.520U
M24     U67_drain D       U48_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.447U PD=.520U
M25     VDD     U43_gate U67_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.520U
M26     VDD     CDN     U48_drain VDD     P   L=0.184U  W=1.91U     
+  PS=.447U
M27     u7_G    E       VSS     VSS     N   L=0.18U  W=0.66U    
M28     u7_G    E       VDD     VDD     P   L=0.18U  W=1.54U    
M29     u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.66U    
M30     u7_GB   u7_G    VDD     VDD     P   L=0.185U  W=1.54U    
M31     U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U    
M32     U43_gate U68_gate VDD     VDD     P   L=0.18U  W=1.8U    
M33     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U    
M34     U68_gate SC      VDD     VDD     P   L=0.184U  W=1.91U    
M35     u9_S    U78_in  VSS     VSS     N   L=0.18U  W=0.83U    
M36     u9_S    U78_in  VDD     VDD     P   L=0.184U  W=1.87U    
M37     U78_in  u9_D    VSS     VSS     N   L=0.18U  W=0.86U    
M38     U78_in  u9_D    VDD     VDD     P   L=0.184U  W=1.87U    
M39     Q       U20_in  VSS     VSS     N   L=0.18U  W=1.38U    
M40     Q       U20_in  VDD     VDD     P   L=0.184U  W=4.1U    
M41     QN      U83_in  VSS     VSS     N   L=0.18U  W=1.38U    
M42     QN      U83_in  VDD     VDD     P   L=0.1845U  W=4.1U    
M43     U83_in  U76_out VSS     VSS     N   L=0.18U  W=0.69U    
M44     U83_in  U76_out VDD     VDD     P   L=0.185U  W=1.76U    
M45     U20_in  U82_out VSS     VSS     N   L=0.18U  W=0.69U    
M46     U20_in  U82_out VDD     VDD     P   L=0.184U  W=2.05U    
M47     SO      U78_in  VSS     VSS     N   L=0.186U  W=1.38U    
M48     SO      U78_in  VDD     VDD     P   L=0.182U  W=4.1U    

.ENDS slbhb2

.SUBCKT slbhb4 SO Q QN  CDN D E SC SD SDN VDD VSS
M1      U82_out SDN     VDD     VDD     P   L=0.184U  W=1.83U    
M2      U82_out U82_in1 VDD     VDD     P   L=0.18U  W=1.83U    
M3      U82_$$7 SDN     VSS     VSS     N   L=0.18U  W=0.83U    
M4      U82_out U82_in1 U82_$$7 VSS     N   L=0.18U  W=0.83U    
M5      U76_out CDN     VDD     VDD     P   L=0.185U  W=1.7U    
M6      U76_out U82_out VDD     VDD     P   L=0.185U  W=1.68U    
M7      U76_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.83U    
M8      U76_out U82_out U76_$$7 VSS     N   L=0.18U  W=0.83U    
M9      U76_out u7_GB   U82_in1 VDD     P   L=0.18U  W=1.41U    
M10     U76_out u7_G    U82_in1 VSS     N   L=0.18U  W=0.46U    
M11     U48_drain u7_G    U82_in1 VDD     P   L=0.185U  W=1.41U     
+  PD=.447U
M12     U48_drain u7_GB   U82_in1 VSS     N   L=0.18U  W=0.46U     
+  PD=.480U
M13     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.82U    
M14     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.54U    
M15     U82_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.82U    
M16     U82_out u7_G    u9_D    VSS     N   L=0.18U  W=0.54U    
M17     U48_drain D       U48_source VSS     N   L=0.18U  W=0.68U     
+  PS=.480U PD=.480U
M18     U48_source U68_gate U68_source VSS     N   L=0.18U  W=0.68U     
+  PS=.420U PD=.480U
M19     U69_drain U43_gate U68_source VSS     N   L=0.18U  W=0.68U     
+  PS=.420U PD=.480U
M20     U68_source CDN     VSS     VSS     N   L=0.18U  W=0.69U     
+  PD=.420U
M21     U48_drain SD      U69_drain VSS     N   L=0.18U  W=0.68U     
+  PS=.480U PD=.480U
M22     U66_drain SD      U48_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.447U PD=.520U
M23     VDD     U68_gate U66_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.520U
M24     U67_drain D       U48_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.447U PD=.520U
M25     VDD     U43_gate U67_drain VDD     P   L=0.18U  W=1.59U     
+  PS=.520U
M26     VDD     CDN     U48_drain VDD     P   L=0.184U  W=1.91U     
+  PS=.447U
M27     u7_G    E       VSS     VSS     N   L=0.18U  W=0.66U    
M28     u7_G    E       VDD     VDD     P   L=0.185U  W=1.54U    
M29     u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.66U    
M30     u7_GB   u7_G    VDD     VDD     P   L=0.18U  W=1.54U    
M31     U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U    
M32     U43_gate U68_gate VDD     VDD     P   L=0.18U  W=1.8U    
M33     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U    
M34     U68_gate SC      VDD     VDD     P   L=0.184U  W=1.91U    
M35     u9_S    U78_in  VSS     VSS     N   L=0.18U  W=0.83U    
M36     u9_S    U78_in  VDD     VDD     P   L=0.184U  W=1.87U    
M37     U78_in  u9_D    VSS     VSS     N   L=0.18U  W=0.86U    
M38     U78_in  u9_D    VDD     VDD     P   L=0.184U  W=1.87U    
M39     Q       U20_in  VSS     VSS     N   L=0.18U  W=2.77U    
M40     Q       U20_in  VDD     VDD     P   L=0.182U  W=8.2U    
M41     QN      U83_in  VSS     VSS     N   L=0.18U  W=2.77U    
M42     QN      U83_in  VDD     VDD     P   L=0.18325U  W=8.2U    
M43     U83_in  U76_out VSS     VSS     N   L=0.18U  W=0.69U    
M44     U83_in  U76_out VDD     VDD     P   L=0.185U  W=1.66U    
M45     U20_in  U82_out VSS     VSS     N   L=0.18U  W=0.69U    
M46     U20_in  U82_out VDD     VDD     P   L=0.184U  W=2.05U    
M47     SO      U78_in  VSS     VSS     N   L=0.18U  W=2.77U    
M48     SO      U78_in  VDD     VDD     P   L=0.182U  W=8.2U    

.ENDS slbhb4

.SUBCKT slchq1 SO Q  CDN D E SC SD VDD VSS
M1      U79_out U79_in  VSS     VSS     N   L=0.18U  W=0.83U  
M2      U79_out U79_in  VDD     VDD     P   L=0.184U  W=1.83U  
M3      SO      u3_in   VSS     VSS     N   L=0.18U  W=0.69U  
M4      SO      u3_in   VDD     VDD     P   L=0.184U  W=2.05U  
M5      u3_in   u8_D    VSS     VSS     N   L=0.18U  W=0.83U  
M6      u3_in   u8_D    VDD     VDD     P   L=0.184U  W=1.88U  
M7      u8_G    E       VSS     VSS     N   L=0.18U  W=0.66U  
M8      u8_G    E       VDD     VDD     P   L=0.185U  W=1.54U  
M9      u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.66U  
M10     u8_GB   u8_G    VDD     VDD     P   L=0.185U  W=1.54U  
M11     U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M12     U43_gate U45_gate VDD     VDD     P   L=0.18U  W=1.8U  
M13     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M14     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M15     U78_out u3_in   VSS     VSS     N   L=0.18U  W=0.83U  
M16     U78_out u3_in   VDD     VDD     P   L=0.184U  W=1.88U  
M17     Q       U79_in  VSS     VSS     N   L=0.18U  W=0.69U  
M18     Q       U79_in  VDD     VDD     P   L=0.184U  W=2.05U  
M19     U76_out CDN     VDD     VDD     P   L=0.18U  W=1.7U  
M20     U76_out U79_out VDD     VDD     P   L=0.185U  W=1.68U  
M21     U76_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.83U  
M22     U76_out U79_out U76_$$7 VSS     N   L=0.18U  W=0.83U  
M23     U79_out u8_GB   u8_D    VDD     P   L=0.18U  W=0.8U  
M24     U79_out u8_G    u8_D    VSS     N   L=0.18U  W=0.46U  
M25     U15_S   u8_G    U79_in  VDD     P   L=0.185U  W=1.41U   PD=.447U
M26     U15_S   u8_GB   U79_in  VSS     N   L=0.18U  W=0.46U   PD=.480U
M27     U76_out u8_GB   U79_in  VDD     P   L=0.18U  W=1.41U  
M28     U76_out u8_G    U79_in  VSS     N   L=0.18U  W=0.46U  
M29     U78_out u8_G    u8_D    VDD     P   L=0.18U  W=0.8U  
M30     U78_out u8_GB   u8_D    VSS     N   L=0.18U  W=0.46U  
M31     VDD     CDN     U15_S   VDD     P   L=0.184U  W=1.91U   PS=.447U
M32     VDD     U43_gate U43_source VDD     P   L=0.186U  W=1.59U   
+  PS=.520U
M33     U43_source D       U15_S   VDD     P   L=0.186U  W=1.59U   
+  PS=.447U PD=.520U
M34     VDD     U45_gate U45_source VDD     P   L=0.18U  W=1.59U   
+  PS=.520U
M35     U45_source SD      U15_S   VDD     P   L=0.18U  W=1.59U   
+  PS=.447U PD=.520U
M36     U68_drain U45_gate U68_source VSS     N   L=0.18U  W=0.68U   
+  PS=.420U PD=.480U
M37     U69_drain U43_gate U68_source VSS     N   L=0.18U  W=0.68U   
+  PS=.420U PD=.480U
M38     U15_S   D       U68_drain VSS     N   L=0.18U  W=0.68U   
+  PS=.480U PD=.480U
M39     U68_source CDN     VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.420U
M40     U15_S   SD      U69_drain VSS     N   L=0.18U  W=0.68U   
+  PS=.480U PD=.480U

.ENDS slchq1

.SUBCKT slchq2 SO Q  CDN D E SC SD VDD VSS
M1      U79_out U79_in  VSS     VSS     N   L=0.18U  W=0.83U  
M2      U79_out U79_in  VDD     VDD     P   L=0.184U  W=1.83U  
M3      SO      u3_in   VSS     VSS     N   L=0.18U  W=1.38U  
M4      SO      u3_in   VDD     VDD     P   L=0.184U  W=4.1U  
M5      u3_in   u8_D    VSS     VSS     N   L=0.18U  W=0.83U  
M6      u3_in   u8_D    VDD     VDD     P   L=0.184U  W=1.88U  
M7      u8_G    E       VSS     VSS     N   L=0.18U  W=0.66U  
M8      u8_G    E       VDD     VDD     P   L=0.185U  W=1.54U  
M9      u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.66U  
M10     u8_GB   u8_G    VDD     VDD     P   L=0.185U  W=1.54U  
M11     U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M12     U43_gate U45_gate VDD     VDD     P   L=0.18U  W=1.8U  
M13     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M14     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M15     U78_out u3_in   VSS     VSS     N   L=0.18U  W=0.83U  
M16     U78_out u3_in   VDD     VDD     P   L=0.184U  W=1.88U  
M17     Q       U79_in  VSS     VSS     N   L=0.18U  W=1.38U  
M18     Q       U79_in  VDD     VDD     P   L=0.184U  W=4.1U  
M19     U76_out CDN     VDD     VDD     P   L=0.18U  W=1.7U  
M20     U76_out U79_out VDD     VDD     P   L=0.185U  W=1.68U  
M21     U76_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.83U  
M22     U76_out U79_out U76_$$7 VSS     N   L=0.18U  W=0.83U  
M23     U79_out u8_GB   u8_D    VDD     P   L=0.18U  W=0.8U  
M24     U79_out u8_G    u8_D    VSS     N   L=0.18U  W=0.46U  
M25     U15_S   u8_G    U79_in  VDD     P   L=0.185U  W=1.41U   PD=.447U
M26     U15_S   u8_GB   U79_in  VSS     N   L=0.18U  W=0.46U   PD=.480U
M27     U76_out u8_GB   U79_in  VDD     P   L=0.18U  W=1.41U  
M28     U76_out u8_G    U79_in  VSS     N   L=0.18U  W=0.46U  
M29     U78_out u8_G    u8_D    VDD     P   L=0.18U  W=0.8U  
M30     U78_out u8_GB   u8_D    VSS     N   L=0.18U  W=0.46U  
M31     VDD     CDN     U15_S   VDD     P   L=0.184U  W=1.91U   PS=.447U
M32     VDD     U43_gate U43_source VDD     P   L=0.186U  W=1.59U   
+  PS=.520U
M33     U43_source D       U15_S   VDD     P   L=0.186U  W=1.59U   
+  PS=.447U PD=.520U
M34     VDD     U45_gate U45_source VDD     P   L=0.18U  W=1.59U   
+  PS=.520U
M35     U45_source SD      U15_S   VDD     P   L=0.18U  W=1.59U   
+  PS=.447U PD=.520U
M36     U68_drain U45_gate U68_source VSS     N   L=0.18U  W=0.68U   
+  PS=.420U PD=.480U
M37     U69_drain U43_gate U68_source VSS     N   L=0.18U  W=0.68U   
+  PS=.420U PD=.480U
M38     U15_S   D       U68_drain VSS     N   L=0.18U  W=0.68U   
+  PS=.480U PD=.480U
M39     U68_source CDN     VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.420U
M40     U15_S   SD      U69_drain VSS     N   L=0.18U  W=0.68U   
+  PS=.480U PD=.480U

.ENDS slchq2

.SUBCKT slchq4 SO Q  CDN D E SC SD VDD VSS
M1      U79_out U79_in  VSS     VSS     N   L=0.18U  W=0.83U  
M2      U79_out U79_in  VDD     VDD     P   L=0.184U  W=1.83U  
M3      SO      u3_in   VSS     VSS     N   L=0.18U  W=2.77U  
M4      SO      u3_in   VDD     VDD     P   L=0.184U  W=8.2U  
M5      u3_in   u8_D    VSS     VSS     N   L=0.18U  W=0.83U  
M6      u3_in   u8_D    VDD     VDD     P   L=0.184U  W=1.88U  
M7      u8_G    E       VSS     VSS     N   L=0.18U  W=0.66U  
M8      u8_G    E       VDD     VDD     P   L=0.185U  W=1.54U  
M9      u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.66U  
M10     u8_GB   u8_G    VDD     VDD     P   L=0.185U  W=1.54U  
M11     U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U  
M12     U43_gate U45_gate VDD     VDD     P   L=0.18U  W=1.8U  
M13     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M14     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M15     U78_out u3_in   VSS     VSS     N   L=0.18U  W=0.83U  
M16     U78_out u3_in   VDD     VDD     P   L=0.184U  W=1.88U  
M17     Q       U79_in  VSS     VSS     N   L=0.18U  W=2.77U  
M18     Q       U79_in  VDD     VDD     P   L=0.183U  W=8.2U  
M19     U76_out CDN     VDD     VDD     P   L=0.18U  W=1.7U  
M20     U76_out U79_out VDD     VDD     P   L=0.185U  W=1.68U  
M21     U76_$$7 CDN     VSS     VSS     N   L=0.18U  W=0.83U  
M22     U76_out U79_out U76_$$7 VSS     N   L=0.18U  W=0.83U  
M23     U79_out u8_GB   u8_D    VDD     P   L=0.18U  W=0.8U  
M24     U79_out u8_G    u8_D    VSS     N   L=0.18U  W=0.46U  
M25     U15_S   u8_G    U79_in  VDD     P   L=0.185U  W=1.41U   PD=.447U
M26     U15_S   u8_GB   U79_in  VSS     N   L=0.18U  W=0.46U   PD=.480U
M27     U76_out u8_GB   U79_in  VDD     P   L=0.18U  W=1.41U  
M28     U76_out u8_G    U79_in  VSS     N   L=0.18U  W=0.46U  
M29     U78_out u8_G    u8_D    VDD     P   L=0.18U  W=0.8U  
M30     U78_out u8_GB   u8_D    VSS     N   L=0.18U  W=0.46U  
M31     VDD     CDN     U15_S   VDD     P   L=0.184U  W=1.91U   PS=.447U
M32     VDD     U43_gate U43_source VDD     P   L=0.186U  W=1.59U   
+  PS=.520U
M33     U43_source D       U15_S   VDD     P   L=0.186U  W=1.59U   
+  PS=.447U PD=.520U
M34     VDD     U45_gate U45_source VDD     P   L=0.18U  W=1.59U   
+  PS=.520U
M35     U45_source SD      U15_S   VDD     P   L=0.18U  W=1.59U   
+  PS=.447U PD=.520U
M36     U68_drain U45_gate U68_source VSS     N   L=0.18U  W=0.68U   
+  PS=.420U PD=.480U
M37     U69_drain U43_gate U68_source VSS     N   L=0.18U  W=0.68U   
+  PS=.420U PD=.480U
M38     U15_S   D       U68_drain VSS     N   L=0.18U  W=0.68U   
+  PS=.480U PD=.480U
M39     U68_source CDN     VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.420U
M40     U15_S   SD      U69_drain VSS     N   L=0.18U  W=0.68U   
+  PS=.480U PD=.480U

.ENDS slchq4

.SUBCKT slclq1 SO Q  CDN D EN SC SD VDD VSS
M1      U79_out U79_in  VSS     VSS     N   L=0.18U  W=0.83U
M2      U79_out U79_in  VDD     VDD     P   L=0.184U  W=1.81U
M3      SO      u3_in   VSS     VSS     N   L=0.18U  W=0.69U
M4      SO      u3_in   VDD     VDD     P   L=0.184U  W=2.05U
M5      u3_in   u8_D    VSS     VSS     N   L=0.18U  W=0.83U
M6      u3_in   u8_D    VDD     VDD     P   L=0.18U  W=1.88U
M7      u8_GB   EN      VSS     VSS     N   L=0.18U  W=0.66U
M8      u8_GB   EN      VDD     VDD     P   L=0.185U  W=1.54U
M9      u8_G    u8_GB   VSS     VSS     N   L=0.18U  W=0.66U
M10     u8_G    u8_GB   VDD     VDD     P   L=0.185U  W=1.54U
M11     U43_gate U45_gate VSS     VSS     N   L=0.18U   W=0.69U
M12     U43_gate U45_gate VDD     VDD     P   L=0.18U   W=1.8U
M13     U45_gate SC      VSS     VSS     N   L=0.18U    W=0.69U
M14     U45_gate SC      VDD     VDD     P   L=0.184U    W=1.91U
M15     U78_out u3_in   VSS     VSS     N   L=0.18U     W=0.83U
M16     U78_out u3_in   VDD     VDD     P   L=0.184U     W=1.88U
M17     Q       U79_in  VSS     VSS     N   L=0.18U     W=0.69U
M18     Q       U79_in  VDD     VDD     P   L=0.184U     W=2.05U
M19     U76_out CDN     VDD     VDD     P   L=0.18U     W=1.70U
M20     U76_out U79_out VDD     VDD     P   L=0.185U     W=1.68U
M21     U76_$$7 CDN     VSS     VSS     N   L=0.18U     W=0.83U
M22     U76_out U79_out U76_$$7 VSS     N   L=0.18U     W=0.83U
M23     U79_out u8_GB   u8_D    VDD     P   L=0.18U     W=0.78U
M24     U79_out u8_G    u8_D    VSS     N   L=0.18U     W=0.46U
M25     U15_S   u8_G    U79_in  VDD     P   L=0.186U     PD=.447U  W=1.34U
M26     U15_S   u8_GB   U79_in  VSS     N   L=0.18U     PD=.480U  W=0.46U
M27     U76_out u8_GB   U79_in  VDD     P   L=0.18U     W=1.38U
M28     U76_out u8_G    U79_in  VSS     N   L=0.18U     W=0.46U
M29     U78_out u8_G    u8_D    VDD     P   L=0.18U     W=0.78U
M30     U78_out u8_GB   u8_D    VSS     N   L=0.18U     W=0.46U
M31     VDD     CDN     U15_S   VDD     P   L=0.184U     PS=.447U  W=1.91U
M32     VDD     U43_gate U43_source VDD     P   L=0.185U      W=1.50U
+  PS=.520U
M33     U43_source D       U15_S   VDD     P   L=0.185U       W=1.50U
+  PS=.447U PD=.520U
M34     VDD     U45_gate U45_source VDD     P   L=0.18U      W=1.59U
+  PS=.520U
M35     U45_source SD      U15_S   VDD     P   L=0.18U       W=1.59U
+  PS=.447U PD=.520U
M36     U68_drain U45_gate U68_source VSS     N   L=0.18U    W=0.68U
+  PS=.420U PD=.480U
M37     U69_drain U43_gate U68_source VSS     N   L=0.18U    W=0.68U
+  PS=.420U PD=.480U
M38     U15_S   D       U68_drain VSS     N   L=0.18U        W=0.68U
+  PS=.480U PD=.480U
M39     U68_source CDN     VSS     VSS     N   L=0.18U       W=0.69U
+  PD=.420U
M40     U15_S   SD      U69_drain VSS     N   L=0.18U        W=0.68U
+  PS=.480U PD=.480U

.ENDS slclq1

.SUBCKT slclq2 SO Q  CDN D EN SC SD VDD VSS
M1      U79_out U79_in  VSS     VSS     N   L=0.18U      W=0.83U
M2      U79_out U79_in  VDD     VDD     P   L=0.184U      W=1.81U
M3      SO      u3_in   VSS     VSS     N   L=0.18U      W=1.38U
M4      SO      u3_in   VDD     VDD     P   L=0.184U      W=4.1U
M5      u3_in   u8_D    VSS     VSS     N   L=0.18U      W=0.83U
M6      u3_in   u8_D    VDD     VDD     P   L=0.18U      W=1.88U
M7      u8_GB   EN      VSS     VSS     N   L=0.18U      W=0.66U
M8      u8_GB   EN      VDD     VDD     P   L=0.185U      W=1.54U
M9      u8_G    u8_GB   VSS     VSS     N   L=0.18U      W=0.66U
M10     u8_G    u8_GB   VDD     VDD     P   L=0.185U      W=1.54U
M11     U43_gate U45_gate VSS     VSS     N   L=0.18U      W=0.69U
M12     U43_gate U45_gate VDD     VDD     P   L=0.18U      W=1.8U
M13     U45_gate SC      VSS     VSS     N   L=0.18U       W=0.69U
M14     U45_gate SC      VDD     VDD     P   L=0.184U       W=1.91U
M15     U78_out u3_in   VSS     VSS     N   L=0.18U        W=0.83U
M16     U78_out u3_in   VDD     VDD     P   L=0.184U        W=1.88U
M17     Q       U79_in  VSS     VSS     N   L=0.18U        W=1.38U
M18     Q       U79_in  VDD     VDD     P   L=0.184U      W=4.1U
M19     U76_out CDN     VDD     VDD     P   L=0.18U      W=1.70U
M20     U76_out U79_out VDD     VDD     P   L=0.185U      W=1.68U
M21     U76_$$7 CDN     VSS     VSS     N   L=0.18U      W=0.83U
M22     U76_out U79_out U76_$$7 VSS     N   L=0.18U      W=0.83U
M23     U79_out u8_GB   u8_D    VDD     P   L=0.18U      W=0.78U
M24     U79_out u8_G    u8_D    VSS     N   L=0.18U      W=0.46U
M25     U15_S   u8_G    U79_in  VDD     P   L=0.186U     PD=.447U  W=1.34U
M26     U15_S   u8_GB   U79_in  VSS     N   L=0.18U     PD=.480U  W=0.46U
M27     U76_out u8_GB   U79_in  VDD     P   L=0.18U      W=1.38U
M28     U76_out u8_G    U79_in  VSS     N   L=0.18U      W=0.46U
M29     U78_out u8_G    u8_D    VDD     P   L=0.18U      W=0.78U
M30     U78_out u8_GB   u8_D    VSS     N   L=0.18U      W=0.46U
M31     VDD     CDN     U15_S   VDD     P   L=0.184U     PS=.447U  W=1.91U
M32     VDD     U43_gate U43_source VDD     P   L=0.185U       W=1.5U
+  PS=.520U
M33     U43_source D       U15_S   VDD     P   L=0.185U       W=1.5U
+  PS=.447U PD=.520U
M34     VDD     U45_gate U45_source VDD     P   L=0.18U       W=1.59U
+  PS=.520U
M35     U45_source SD      U15_S   VDD     P   L=0.18U       W=1.59U
+  PS=.447U PD=.520U
M36     U68_drain U45_gate U68_source VSS     N   L=0.18U       W=0.68U
+  PS=.420U PD=.480U
M37     U69_drain U43_gate U68_source VSS     N   L=0.18U       W=0.68U
+  PS=.420U PD=.480U
M38     U15_S   D       U68_drain VSS     N   L=0.18U       W=0.68U
+  PS=.480U PD=.480U
M39     U68_source CDN     VSS     VSS     N   L=0.18U       W=0.69U
+  PD=.420U
M40     U15_S   SD      U69_drain VSS     N   L=0.18U       W=0.68U
+  PS=.480U PD=.480U

.ENDS slclq2

.SUBCKT slclq4 SO Q  CDN D EN SC SD VDD VSS
M1      U79_out U79_in  VSS     VSS     N   L=0.18U      W=0.83U
M2      U79_out U79_in  VDD     VDD     P   L=0.184U      W=1.81U
M3      SO      u3_in   VSS     VSS     N   L=0.18U      W=2.77U
M4      SO      u3_in   VDD     VDD     P   L=0.184U      W=8.2U
M5      u3_in   u8_D    VSS     VSS     N   L=0.18U      W=0.83U
M6      u3_in   u8_D    VDD     VDD     P   L=0.18U      W=1.89U
M7      u8_GB   EN      VSS     VSS     N   L=0.18U      W=0.66U
M8      u8_GB   EN      VDD     VDD     P   L=0.185U      W=1.54U
M9      u8_G    u8_GB   VSS     VSS     N   L=0.18U      W=0.66U
M10     u8_G    u8_GB   VDD     VDD     P   L=0.185U      W=1.54U
M11     U43_gate U45_gate VSS     VSS     N   L=0.18U      W=0.69U
M12     U43_gate U45_gate VDD     VDD     P   L=0.18U      W=1.8U
M13     U45_gate SC      VSS     VSS     N   L=0.18U      W=0.69U
M14     U45_gate SC      VDD     VDD     P   L=0.184U      W=1.91U
M15     U78_out u3_in   VSS     VSS     N   L=0.18U      W=0.83U
M16     U78_out u3_in   VDD     VDD     P   L=0.184U      W=1.89U
M17     Q       U79_in  VSS     VSS     N   L=0.18U     W=2.77U
M18     Q       U79_in  VDD     VDD     P   L=0.183U      W=8.2U
M19     U76_out CDN     VDD     VDD     P   L=0.18U      W=1.70U
M20     U76_out U79_out VDD     VDD     P   L=0.185U      W=1.68U
M21     U76_$$7 CDN     VSS     VSS     N   L=0.18U      W=0.83U
M22     U76_out U79_out U76_$$7 VSS     N   L=0.18U      W=0.83U
M23     U79_out u8_GB   u8_D    VDD     P   L=0.18U      W=0.78U
M24     U79_out u8_G    u8_D    VSS     N   L=0.18U      W=0.46U
M25     U15_S   u8_G    U79_in  VDD     P   L=0.186U     PD=.447U  W=1.34U
M26     U15_S   u8_GB   U79_in  VSS     N   L=0.18U     PD=.480U  W=0.46U
M27     U76_out u8_GB   U79_in  VDD     P   L=0.18U      W=1.38U
M28     U76_out u8_G    U79_in  VSS     N   L=0.18U      W=0.46U
M29     U78_out u8_G    u8_D    VDD     P   L=0.18U      W=0.78U
M30     U78_out u8_GB   u8_D    VSS     N   L=0.18U      W=0.46U
M31     VDD     CDN     U15_S   VDD     P   L=0.184U     PS=.447U  W=1.91U
M32     VDD     U43_gate U43_source VDD     P   L=0.185U       W=1.50U
+  PS=.520U
M33     U43_source D       U15_S   VDD     P   L=0.185U       W=1.50U
+  PS=.447U PD=.520U
M34     VDD     U45_gate U45_source VDD     P   L=0.18U       W=1.59U
+  PS=.520U
M35     U45_source SD      U15_S   VDD     P   L=0.18U       W=1.59U
+  PS=.447U PD=.520U
M36     U68_drain U45_gate U68_source VSS     N   L=0.18U       W=0.68U
+  PS=.420U PD=.480U
M37     U69_drain U43_gate U68_source VSS     N   L=0.18U       W=0.68U
+  PS=.420U PD=.480U
M38     U15_S   D       U68_drain VSS     N   L=0.18U       W=0.68U
+  PS=.480U PD=.480U
M39     U68_source CDN     VSS     VSS     N   L=0.18U       W=0.69U
+  PD=.420U
M40     U15_S   SD      U69_drain VSS     N   L=0.18U       W=0.68U
+  PS=.480U PD=.480U

.ENDS slclq4

.SUBCKT slnhb1 SO Q QN  D E SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.83U
M2      U35_out U35_in  VDD     VDD     P   L=0.18U  W=1.83U
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.83U
M4      U37_out U35_out VDD     VDD     P   L=0.18U  W=1.83U
M5      SO      u3_in   VSS     VSS     N   L=0.18U  W=0.69U
M6      SO      u3_in   VDD     VDD     P   L=0.184U W=2.05U
M7      u3_in   U38_in  VSS     VSS     N   L=0.18U  W=0.83U
M8      u3_in   U38_in  VDD     VDD     P   L=0.185U  W=1.805U
M9      u8_G    E       VSS     VSS     N   L=0.18U  W=0.66U
M10     u8_G    E       VDD     VDD     P   L=0.184U  W=1.74U
M11     u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.66U
M12     u8_GB   u8_G    VDD     VDD     P   L=0.184U  W=1.74U
M13     U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U
M14     U43_gate U45_gate VDD     VDD     P   L=0.18U  W=1.91U
M15     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U
M16     U45_gate SC      VDD     VDD     P   L=0.184U W=1.91U
M17     U36_out u3_in   VSS     VSS     N   L=0.18U  W=0.83U
M18     U36_out u3_in   VDD     VDD     P   L=0.185U  W=1.805U
M19     QN      U35_out VSS     VSS     N   L=0.18U  W=0.69U
M20     QN      U35_out VDD     VDD     P   L=0.185U  W=1.977U
M21     Q       U35_in  VSS     VSS     N   L=0.18U  W=0.69U
M22     Q       U35_in  VDD     VDD     P   L=0.187U  W=1.954U
M23     U35_out u8_GB   U38_in  VDD     P   L=0.18U  W=0.69U
M24     U35_out u8_G    U38_in  VSS     N   L=0.18U  W=0.46U
M25     U15_S   u8_G    U35_in  VDD     P   L=0.18U  W=1.44U
M26     U15_S   u8_GB   U35_in  VSS     N   L=0.18U  W=0.46U
M27     U37_out u8_GB   U35_in  VDD     P   L=0.186U  W=1.44U
M28     U37_out u8_G    U35_in  VSS     N   L=0.18U  W=0.46U
M29     U36_out u8_G    U38_in  VDD     P   L=0.18U  W=0.69U
M30     U36_out u8_GB   U38_in  VSS     N   L=0.18U  W=0.42U
M31     VDD     U45_gate U45_source VDD     P   L=0.18U  W=1.91U
+  PS=.520U
M32     U45_source SD      U15_S   VDD     P   L=0.18U  W=1.91U
+  PS=.520U PD=.520U
M33     U67_drain D       U15_S   VDD     P   L=0.185U  W=1.78U
+  PS=.520U PD=.520U
M34     VDD     U43_gate U67_drain VDD     P   L=0.185U  W=1.78U
+  PS=.520U
M35     U15_S   D       U48_source VSS     N   L=0.18U  W=0.69U
+  PS=.480U PD=.480U
M36     U48_source U45_gate VSS     VSS     N   L=0.18U  W=0.69U
+  PD=.480U
M37     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U
+  PD=.480U
M38     U15_S   SD      U69_drain VSS     N   L=0.18U  W=0.66U
+  PS=.480U PD=.480U

.ENDS slnhb1

.SUBCKT slnhb2 SO Q QN  D E SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.83U
M2      U35_out U35_in  VDD     VDD     P   L=0.18U  W=1.83U
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.83U
M4      U37_out U35_out VDD     VDD     P   L=0.18U  W=1.83U
M5      SO      u3_in   VSS     VSS     N   L=0.18U  W=1.38U
M6      SO      u3_in   VDD     VDD     P   L=0.1875U  W=4.1U
M7      u3_in   U38_in  VSS     VSS     N   L=0.18U  W=0.83U
M8      u3_in   U38_in  VDD     VDD     P   L=0.18U  W=1.88U
M9      u8_G    E       VSS     VSS     N   L=0.18U  W=0.66U
M10     u8_G    E       VDD     VDD     P   L=0.184U  W=1.74U
M11     u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.66U
M12     u8_GB   u8_G    VDD     VDD     P   L=0.18U  W=1.74U
M13     U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U
M14     U43_gate U68_gate VDD     VDD     P   L=0.18U  W=1.91U
M15     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U
M16     U68_gate SC      VDD     VDD     P   L=0.184U  W=1.91U
M17     u9_S    u3_in   VSS     VSS     N   L=0.18U  W=0.83U
M18     u9_S    u3_in   VDD     VDD     P   L=0.184U  W=1.88U
M19     Q       U35_in  VSS     VSS     N   L=0.18U  W=1.38U
M20     Q       U35_in  VDD     VDD     P   L=0.186U  W=4.1U
M21     QN      U35_out VSS     VSS     N   L=0.18U  W=1.38U
M22     QN      U35_out VDD     VDD     P   L=0.1865U  W=4.1U
M23     VDD     U43_gate U43_source VDD     P   L=0.185U  W=1.78U
+  PS=.520U
M24     U43_source D       U67_source VDD     P   L=0.185U  W=1.78U
+  PS=.520U PD=.520U
M25     VDD     U68_gate U45_source VDD     P   L=0.18U  W=1.91U
+  PS=.520U
M26     U45_source SD      U67_source VDD     P   L=0.18U  W=1.91U
+  PS=.520U PD=.520U
M27     U68_drain U68_gate VSS     VSS     N   L=0.18U  W=0.69U
+  PD=.480U
M28     U67_source D       U68_drain VSS     N   L=0.18U  W=0.69U
+  PS=.480U PD=.480U
M29     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U
+  PD=.480U
M30     U67_source SD      U69_drain VSS     N   L=0.18U  W=0.66U
+  PS=.480U PD=.480U
M31     U35_out u8_GB   U38_in  VDD     P   L=0.18U  W=0.69U
M32     U35_out u8_G    U38_in  VSS     N   L=0.18U  W=0.46U
M33     U67_source u8_G    U35_in  VDD     P   L=0.18U  W=1.44U
+  PD=.520U
M34     U67_source u8_GB   U35_in  VSS     N   L=0.18U  W=0.46U
+  PD=.480U
M35     U37_out u8_GB   U35_in  VDD     P   L=0.186U  W=1.44U
M36     U37_out u8_G    U35_in  VSS     N   L=0.18U  W=0.46U
M37     u9_S    u8_G    U38_in  VDD     P   L=0.18U  W=0.69U
M38     u9_S    u8_GB   U38_in  VSS     N   L=0.18U  W=0.42U

.ENDS slnhb2

.SUBCKT slnhb4 SO Q QN  D E SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.83U
M2      U35_out U35_in  VDD     VDD     P   L=0.18U  W=1.83U
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.83U
M4      U37_out U35_out VDD     VDD     P   L=0.184U  W=1.83U
M5      SO      u3_in   VSS     VSS     N   L=0.18U  W=2.77U
M6      SO      u3_in   VDD     VDD     P   L=0.18725U  W=8.2U
M7      u3_in   U38_in  VSS     VSS     N   L=0.18U  W=0.83U
M8      u3_in   U38_in  VDD     VDD     P   L=0.18U  W=1.88U
M9      u8_G    E       VSS     VSS     N   L=0.18U  W=0.66U
M10     u8_G    E       VDD     VDD     P   L=0.184U  W=1.74U
M11     u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.66U
M12     u8_GB   u8_G    VDD     VDD     P   L=0.184U  W=1.74U
M13     U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U
M14     U43_gate U68_gate VDD     VDD     P   L=0.18U  W=1.91U
M15     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U
M16     U68_gate SC      VDD     VDD     P   L=0.184U  W=1.91U
M17     u9_S    u3_in   VSS     VSS     N   L=0.18U  W=0.83U
M18     u9_S    u3_in   VDD     VDD     P   L=0.184U  W=1.88U
M19     Q       U35_in  VSS     VSS     N   L=0.18U  W=2.77U
M20     Q       U35_in  VDD     VDD     P   L=0.187U  W=8.2U
M21     QN      U35_out VSS     VSS     N   L=0.18U  W=2.77U
M22     QN      U35_out VDD     VDD     P   L=0.187U  W=8.2U
M23     VDD     U43_gate U43_source VDD     P   L=0.185U  W=1.78U
+  PS=.520U
M24     U43_source D       U67_source VDD     P   L=0.185U  W=1.78U
+  PS=.520U PD=.520U
M25     VDD     U68_gate U45_source VDD     P   L=0.18U  W=1.91U
+  PS=.520U
M26     U45_source SD      U67_source VDD     P   L=0.18U  W=1.91U
+  PS=.520U PD=.520U
M27     U68_drain U68_gate VSS     VSS     N   L=0.18U  W=0.69U
+  PD=.480U
M28     U67_source D       U68_drain VSS     N   L=0.18U  W=0.69U
+  PS=.480U PD=.480U
M29     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U
+  PD=.480U
M30     U67_source SD      U69_drain VSS     N   L=0.18U  W=0.66U
+  PS=.480U PD=.480U
M31     U35_out u8_GB   U38_in  VDD     P   L=0.18U  W=0.69U
M32     U35_out u8_G    U38_in  VSS     N   L=0.18U  W=0.46U
M33     U67_source u8_G    U35_in  VDD     P   L=0.18U  W=1.44U
+  PD=.520U
M34     U67_source u8_GB   U35_in  VSS     N   L=0.18U  W=0.46U
+  PD=.480U
M35     U37_out u8_GB   U35_in  VDD     P   L=0.186U  W=1.44U
M36     U37_out u8_G    U35_in  VSS     N   L=0.18U  W=0.46U
M37     u9_S    u8_G    U38_in  VDD     P   L=0.18U  W=0.69U
M38     u9_S    u8_GB   U38_in  VSS     N   L=0.18U  W=0.42U

.ENDS slnhb4

.SUBCKT slnhn1 SO QN  D E SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.83U  
M2      U35_out U35_in  VDD     VDD     P   L=0.184U  W=1.83U  
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.83U  
M4      U37_out U35_out VDD     VDD     P   L=0.18U  W=1.83U  
M5      u7_G    E       VSS     VSS     N   L=0.18U  W=0.66U  
M6      u7_G    E       VDD     VDD     P   L=0.184U  W=1.74U  
M7      u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.66U  
M8      u7_GB   u7_G    VDD     VDD     P   L=0.18U  W=1.74U  
M9      U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U  
M10     U43_gate U68_gate VDD     VDD     P   L=0.184U  W=1.91U  
M11     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M12     U68_gate SC      VDD     VDD     P   L=0.18U  W=1.91U  
M13     u9_S    U36_in  VSS     VSS     N   L=0.18U  W=.83U  
M14     u9_S    U36_in  VDD     VDD     P   L=0.184U  W=1.88U  
M15     QN      U35_out VSS     VSS     N   L=0.18U  W=0.69U  
M16     QN      U35_out VDD     VDD     P   L=0.183U  W=2.05U  
M17     SO      U36_in  VSS     VSS     N   L=0.18U  W=0.69U  
M18     SO      U36_in  VDD     VDD     P   L=0.184U  W=2.05U  
M19     U36_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M20     U36_in  u9_D    VDD     VDD     P   L=0.184U  W=1.88U  
M21     VDD     U43_gate U43_source VDD     P   L=0.184U  W=1.78U   
+  PS=.520U
M22     U43_source D       U67_source VDD     P   L=0.184U  W=1.78U   
+  PS=.520U PD=.520U
M23     VDD     U68_gate U45_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M24     U45_source SD      U67_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M25     U68_drain U68_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M26     U67_source D       U68_drain VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M27     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M28     U67_source SD      U69_drain VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U
M29     U37_out u7_GB   U35_in  VDD     P   L=0.185U  W=1.44U  
M30     U37_out u7_G    U35_in  VSS     N   L=0.18U  W=0.46U  
M31     U67_source u7_G    U35_in  VDD     P   L=0.185U  W=1.44U   
+  PD=.520U
M32     U67_source u7_GB   U35_in  VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M33     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.69U  
M34     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M35     U35_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.69U  
M36     U35_out u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  

.ENDS slnhn1

.SUBCKT slnhn2 SO QN  D E SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.83U  
M2      U35_out U35_in  VDD     VDD     P   L=0.184U  W=1.83U  
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.83U  
M4      U37_out U35_out VDD     VDD     P   L=0.18U  W=1.83U  
M5      u7_G    E       VSS     VSS     N   L=0.18U  W=0.66U  
M6      u7_G    E       VDD     VDD     P   L=0.184U  W=1.74U  
M7      u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.66U  
M8      u7_GB   u7_G    VDD     VDD     P   L=0.18U  W=1.74U  
M9      U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U  
M10     U43_gate U68_gate VDD     VDD     P   L=0.184U  W=1.91U  
M11     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M12     U68_gate SC      VDD     VDD     P   L=0.18U  W=1.91U  
M13     u9_S    U36_in  VSS     VSS     N   L=0.18U  W=.83U  
M14     u9_S    U36_in  VDD     VDD     P   L=0.184U  W=1.88U  
M15     QN      U35_out VSS     VSS     N   L=0.18U  W=1.38U  
M16     QN      U35_out VDD     VDD     P   L=0.183U  W=4.1U  
M17     SO      U36_in  VSS     VSS     N   L=0.18U  W=1.38U  
M18     SO      U36_in  VDD     VDD     P   L=0.183U  W=4.1U  
M19     U36_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M20     U36_in  u9_D    VDD     VDD     P   L=0.18U  W=1.88U  
M21     VDD     U43_gate U43_source VDD     P   L=0.184U  W=1.78U   
+  PS=.520U
M22     U43_source D       U67_source VDD     P   L=0.184U  W=1.78U   
+  PS=.520U PD=.520U
M23     VDD     U68_gate U45_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M24     U45_source SD      U67_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M25     U68_drain U68_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M26     U67_source D       U68_drain VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M27     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M28     U67_source SD      U69_drain VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U
M29     U37_out u7_GB   U35_in  VDD     P   L=0.185U  W=1.44U  
M30     U37_out u7_G    U35_in  VSS     N   L=0.18U  W=0.46U  
M31     U67_source u7_G    U35_in  VDD     P   L=0.185U  W=1.44U   
+  PD=.520U
M32     U67_source u7_GB   U35_in  VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M33     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.69U  
M34     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M35     U35_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.69U  
M36     U35_out u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  

.ENDS slnhn2

.SUBCKT slnhn4 SO QN  D E SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.83U  
M2      U35_out U35_in  VDD     VDD     P   L=0.184U  W=1.83U  
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.83U  
M4      U37_out U35_out VDD     VDD     P   L=0.18U  W=1.83U  
M5      u7_G    E       VSS     VSS     N   L=0.18U  W=0.66U  
M6      u7_G    E       VDD     VDD     P   L=0.184U  W=1.74U  
M7      u7_GB   u7_G    VSS     VSS     N   L=0.18U  W=0.66U  
M8      u7_GB   u7_G    VDD     VDD     P   L=0.18U  W=1.74U  
M9      U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U  
M10     U43_gate U68_gate VDD     VDD     P   L=0.184U  W=1.91U  
M11     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M12     U68_gate SC      VDD     VDD     P   L=0.18U  W=1.91U  
M13     u9_S    U36_in  VSS     VSS     N   L=0.18U  W=.83U  
M14     u9_S    U36_in  VDD     VDD     P   L=0.184U  W=1.88U  
M15     QN      U35_out VSS     VSS     N   L=0.18U  W=2.77U  
M16     QN      U35_out VDD     VDD     P   L=0.183U  W=8.2U  
M17     SO      U36_in  VSS     VSS     N   L=0.18U  W=2.77U  
M18     SO      U36_in  VDD     VDD     P   L=0.183U  W=8.2U  
M19     U36_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M20     U36_in  u9_D    VDD     VDD     P   L=0.18U  W=1.88U  
M21     VDD     U43_gate U43_source VDD     P   L=0.184U  W=1.78U   
+  PS=.520U
M22     U43_source D       U67_source VDD     P   L=0.184U  W=1.78U   
+  PS=.520U PD=.520U
M23     VDD     U68_gate U45_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M24     U45_source SD      U67_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M25     U68_drain U68_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M26     U67_source D       U68_drain VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M27     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M28     U67_source SD      U69_drain VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U
M29     U37_out u7_GB   U35_in  VDD     P   L=0.185U  W=1.44U  
M30     U37_out u7_G    U35_in  VSS     N   L=0.18U  W=0.46U  
M31     U67_source u7_G    U35_in  VDD     P   L=0.185U  W=1.44U   
+  PD=.520U
M32     U67_source u7_GB   U35_in  VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M33     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.69U  
M34     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M35     U35_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.69U  
M36     U35_out u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  

.ENDS slnhn4

.SUBCKT slnhq1 SO Q  D E SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.83U
M2      U35_out U35_in  VDD     VDD     P   L=0.18U  W=1.83U
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.83U
M4      U37_out U35_out VDD     VDD     P   L=0.184U  W=1.83U
M5      SO      u3_in   VSS     VSS     N   L=0.18U  W=0.69U
M6      SO      u3_in   VDD     VDD     P   L=0.184U  W=2.05U
M7      u3_in   u8_D    VSS     VSS     N   L=0.18U  W=0.83U
M8      u3_in   u8_D    VDD     VDD     P   L=0.185U  W=1.88U
M9      u8_G    E       VSS     VSS     N   L=0.18U  W=0.66U
M10     u8_G    E       VDD     VDD     P   L=0.184U  W=1.74U
M11     u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.66U
M12     u8_GB   u8_G    VDD     VDD     P   L=0.184U  W=1.74U
M13     U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U
M14     U43_gate U45_gate VDD     VDD     P   L=0.18U  W=1.91U
M15     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U
M16     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U
M17     U36_out u3_in   VSS     VSS     N   L=0.18U  W=0.83U
M18     U36_out u3_in   VDD     VDD     P   L=0.185U  W=1.792U
M19     Q       U35_in  VSS     VSS     N   L=0.18U  W=0.69U
M20     Q       U35_in  VDD     VDD     P   L=0.1825U  W=2.05U
M21     U35_out u8_GB   u8_D    VDD     P   L=0.18U  W=0.69U
M22     U35_out u8_G    u8_D    VSS     N   L=0.18U  W=0.46U
M23     U15_S   u8_G    U35_in  VDD     P   L=0.18U  W=1.38U
M24     U15_S   u8_GB   U35_in  VSS     N   L=0.18U  W=0.46U
M25     U37_out u8_GB   U35_in  VDD     P   L=0.186U  W=1.38U
M26     U37_out u8_G    U35_in  VSS     N   L=0.18U  W=0.46U
M27     U36_out u8_G    u8_D    VDD     P   L=0.18U  W=0.69U
M28     U36_out u8_GB   u8_D    VSS     N   L=0.18U  W=0.42U
M29     VDD     U45_gate U45_source VDD     P   L=0.18U  W=1.91U
+  PS=.520U
M30     U45_source SD      U15_S   VDD     P   L=0.18U  W=1.91U
+  PS=.520U PD=.520U
M31     U67_drain D       U15_S   VDD     P   L=0.185U  W=1.78U
+  PS=.520U PD=.520U
M32     VDD     U43_gate U67_drain VDD     P   L=0.185U  W=1.78U
+  PS=.520U
M33     U15_S   D       U48_source VSS     N   L=0.18U  W=0.69U
+  PS=.480U PD=.480U
M34     U48_source U45_gate VSS     VSS     N   L=0.18U  W=0.69U
+  PD=.480U
M35     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U
+  PD=.480U
M36     U15_S   SD      U69_drain VSS     N   L=0.18U  W=0.66U
+  PS=.480U PD=.480U

.ENDS slnhq1

.SUBCKT slnhq2 SO Q  D E SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.83U
M2      U35_out U35_in  VDD     VDD     P   L=0.18U  W=1.83U
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.83U
M4      U37_out U35_out VDD     VDD     P   L=0.185U  W=1.83U
M5      SO      u3_in   VSS     VSS     N   L=0.18U  W=1.38U
M6      SO      u3_in   VDD     VDD     P   L=0.1845U  W=3.954U
M7      u3_in   u8_D    VSS     VSS     N   L=0.18U  W=0.83U
M8      u3_in   u8_D    VDD     VDD     P   L=0.18U  W=1.88U
M9      u8_G    E       VSS     VSS     N   L=0.18U  W=0.66U
M10     u8_G    E       VDD     VDD     P   L=0.18U  W=1.74U
M11     u8_GB   u8_G    VSS     VSS     N   L=0.18U  W=0.66U
M12     u8_GB   u8_G    VDD     VDD     P   L=0.18U  W=1.74U
M13     U43_gate U45_gate VSS     VSS     N   L=0.18U  W=0.69U
M14     U43_gate U45_gate VDD     VDD     P   L=0.18U  W=1.91U
M15     U45_gate SC      VSS     VSS     N   L=0.18U  W=0.69U
M16     U45_gate SC      VDD     VDD     P   L=0.184U  W=1.91U
M17     U36_out u3_in   VSS     VSS     N   L=0.18U  W=0.83U
M18     U36_out u3_in   VDD     VDD     P   L=0.185U  W=1.88U
M19     Q       U35_in  VSS     VSS     N   L=0.18U  W=1.38U
M20     Q       U35_in  VDD     VDD     P   L=0.1845U  W=3.954U
M21     U35_out u8_GB   u8_D    VDD     P   L=0.18U  W=0.69U
M22     U35_out u8_G    u8_D    VSS     N   L=0.18U  W=0.46U
M23     U15_S   u8_G    U35_in  VDD     P   L=0.18U  W=1.38U
M24     U15_S   u8_GB   U35_in  VSS     N   L=0.18U  W=0.46U
M25     U37_out u8_GB   U35_in  VDD     P   L=0.186U  W=1.38U
M26     U37_out u8_G    U35_in  VSS     N   L=0.18U  W=0.46U
M27     U36_out u8_G    u8_D    VDD     P   L=0.18U  W=0.69U
M28     U36_out u8_GB   u8_D    VSS     N   L=0.18U  W=0.42U
M29     VDD     U45_gate U45_source VDD     P   L=0.18U  W=1.91U
+  PS=.520U
M30     U45_source SD      U15_S   VDD     P   L=0.18U  W=1.91U
+  PS=.520U PD=.520U
M31     U67_drain D       U15_S   VDD     P   L=0.185U  W=1.78U
+  PS=.520U PD=.520U
M32     VDD     U43_gate U67_drain VDD     P   L=0.185U  W=1.78U
+  PS=.520U
M33     U15_S   D       U48_source VSS     N   L=0.18U  W=0.69U
+  PS=.480U PD=.480U
M34     U48_source U45_gate VSS     VSS     N   L=0.18U  W=0.69U
+  PD=.480U
M35     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U
+  PD=.480U
M36     U15_S   SD      U69_drain VSS     N   L=0.18U  W=0.66U
+  PS=.480U PD=.480U

.ENDS slnhq2

.SUBCKT slnhq4 SO Q  D E SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U      W=0.83U
M2      U35_out U35_in  VDD     VDD     P   L=0.184U      W=1.83U
M3      U37_out U35_out VSS     VSS     N   L=0.18U      W=0.83U
M4      U37_out U35_out VDD     VDD     P   L=0.184U      W=1.83U
M5      SO      u3_in   VSS     VSS     N   L=0.18U      W=2.77U
M6      SO      u3_in   VDD     VDD     P   L=0.183U      W=7.93U
M7      u3_in   u8_D    VSS     VSS     N   L=0.18U      W=0.83U
M8      u3_in   u8_D    VDD     VDD     P   L=0.18U      W=1.88U
M9      u8_G    E       VSS     VSS     N   L=0.18U      W=0.66U
M10     u8_G    E       VDD     VDD     P   L=0.18U      W=1.74U
M11     u8_GB   u8_G    VSS     VSS     N   L=0.18U      W=0.66U
M12     u8_GB   u8_G    VDD     VDD     P   L=0.18U      W=1.74U
M13     U43_gate U45_gate VSS     VSS     N   L=0.18U      W=0.69U
M14     U43_gate U45_gate VDD     VDD     P   L=0.18U      W=1.91U
M15     U45_gate SC      VSS     VSS     N   L=0.18U      W=0.69U
M16     U45_gate SC      VDD     VDD     P   L=0.184U      W=1.91U
M17     U36_out u3_in   VSS     VSS     N   L=0.18U      W=0.83U
M18     U36_out u3_in   VDD     VDD     P   L=0.184U      W=1.87U
M19     Q       U35_in  VSS     VSS     N   L=0.18U      W=2.77U
M20     Q       U35_in  VDD     VDD     P   L=0.183U      W=7.93U
M21     U35_out u8_GB   u8_D    VDD     P   L=0.18U      W=0.69U
M22     U35_out u8_G    u8_D    VSS     N   L=0.18U      W=0.46U
M23     U15_S   u8_G    U35_in  VDD     P   L=0.18U     PD=.520U  W=1.38U
M24     U15_S   u8_GB   U35_in  VSS     N   L=0.18U     PD=.480U  W=0.46U
M25     U37_out u8_GB   U35_in  VDD     P   L=0.186U      W=1.38U
M26     U37_out u8_G    U35_in  VSS     N   L=0.18U      W=0.46U
M27     U36_out u8_G    u8_D    VDD     P   L=0.18U      W=0.69U
M28     U36_out u8_GB   u8_D    VSS     N   L=0.18U      W=0.42U
M29     VDD     U45_gate U45_source VDD     P   L=0.18U       W=1.91U
+  PS=.520U
M30     U45_source SD      U15_S   VDD     P   L=0.18U       W=1.91U
+  PS=.520U PD=.520U
M31     U67_drain D       U15_S   VDD     P   L=0.185U       W=1.78U
+  PS=.520U PD=.520U
M32     VDD     U43_gate U67_drain VDD     P   L=0.185U       W=1.78U
+  PS=.520U
M33     U15_S   D       U48_source VSS     N   L=0.18U       W=0.69U
+  PS=.480U PD=.480U
M34     U48_source U45_gate VSS     VSS     N   L=0.18U       W=0.69U
+  PD=.480U
M35     U69_drain U43_gate VSS     VSS     N   L=0.18U       W=0.66U
+  PD=.480U
M36     U15_S   SD      U69_drain VSS     N   L=0.18U       W=0.66U
+  PS=.480U PD=.480U

.ENDS slnhq4

.SUBCKT slnht1 SO Z  D E OE SC SD VDD VSS
M1      U1_out  OE      VSS     VSS     N   L=0.18U  W=0.69U  
M2      U1_out  OE      VDD     VDD     P   L=0.184U  W=2.04U  
M3      U35_out nint  VSS     VSS     N   L=0.18U  W=0.83U  
M4      U35_out nint  VDD     VDD     P   L=0.18U  W=1.83U  
M5      U72_out SC      VSS     VSS     N   L=0.18U  W=0.69U  
M6      U72_out SC      VDD     VDD     P   L=0.184U  W=1.91U  
M7      U71_out U72_out VSS     VSS     N   L=0.18U  W=0.69U  
M8      U71_out U72_out VDD     VDD     P   L=0.184U  W=1.91U  
M9      u10_out E       VSS     VSS     N   L=0.18U  W=0.66U  
M10     u10_out E       VDD     VDD     P   L=0.184U  W=1.74U  
M11     u11_out u10_out VSS     VSS     N   L=0.18U  W=0.66U  
M12     u11_out u10_out VDD     VDD     P   L=0.184U  W=1.74U  
M13     u7_S    U35_out VSS     VSS     N   L=0.18U  W=0.83U  
M14     u7_S    U35_out VDD     VDD     P   L=0.184U  W=1.83U  
M15     SO      u3_in   VSS     VSS     N   L=0.18U  W=0.69U  
M16     SO      u3_in   VDD     VDD     P   L=0.184U  W=2.05U  
M17     u3_in   u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M18     u3_in   u9_D    VDD     VDD     P   L=0.184U  W=1.88U  
M19     u9_S    u3_in   VSS     VSS     N   L=0.18U  W=.83U  
M20     u9_S    u3_in   VDD     VDD     P   L=0.185U  W=1.88U  
M21     U50_drain SD      U50_source VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U
M22     U50_drain D       U48_source VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M23     U50_source U71_out VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M24     U48_source U72_out VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M25     Z       OE      U53_source VSS     N   L=0.18U  W=0.69U   
+  PS=1.469U PD=1.234U
M26     U53_source nint  VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=1.469U
M27     U6_drain nint  VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=1.000U
M28     Z       OE      U6_drain VSS     N   L=0.18U  W=0.69U   
+  PS=1.000U PD=1.234U
M29     U66_drain SD      U50_drain VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M30     U67_drain D       U50_drain VDD     P   L=0.185U  W=1.78U   
+  PS=.520U PD=.520U
M31     VDD     U71_out U67_drain VDD     P   L=0.185U  W=1.78U   
+  PS=.520U
M32     VDD     U72_out U66_drain VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M33     Z       U1_out  U42_source VDD     P   L=0.18U  W=2.04U   
+  PS=1.613U PD=1.556U
M34     U76_drain nint  VDD     VDD     P   L=0.182U  W=2.04U   
+  PD=1.500U
M35     Z       U1_out  U76_drain VDD     P   L=0.182U  W=2.04U   
+  PS=1.500U PD=1.556U
M36     U42_source nint  VDD     VDD     P   L=0.18U  W=2.04U   
+  PD=1.613U
M37     U50_drain u10_out nint  VDD     P   L=0.18U  W=1.38U   
+  PD=.520U
M38     U50_drain u11_out nint  VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M39     u7_S    u11_out nint  VDD     P   L=0.18U  W=1.38U  
M40     u7_S    u10_out nint  VSS     N   L=0.18U  W=0.46U  
M41     u9_S    u10_out u9_D    VDD     P   L=0.18U  W=0.69U  
M42     u9_S    u11_out u9_D    VSS     N   L=0.18U  W=0.42U  
M43     U35_out u11_out u9_D    VDD     P   L=0.18U  W=0.69U  
M44     U35_out u10_out u9_D    VSS     N   L=0.18U  W=0.46U  

.ENDS slnht1

.SUBCKT slnht2 SO Z  D E OE SC SD VDD VSS
M1      U1_out  OE      VSS     VSS     N   L=0.18U  W=0.69U  
M2      U1_out  OE      VDD     VDD     P   L=0.184U  W=2.05U  
M3      U72_out SC      VSS     VSS     N   L=0.18U  W=0.69U  
M4      U72_out SC      VDD     VDD     P   L=0.184U  W=1.91U  
M5      U71_out U72_out VSS     VSS     N   L=0.18U  W=0.69U  
M6      U71_out U72_out VDD     VDD     P   L=0.184U  W=1.91U  
M7      u10_out E       VSS     VSS     N   L=0.18U  W=0.66U  
M8      u10_out E       VDD     VDD     P   L=0.184U  W=1.74U  
M9      u11_out u10_out VSS     VSS     N   L=0.18U  W=0.66U  
M10     u11_out u10_out VDD     VDD     P   L=0.184U  W=1.74U  
M11     U35_out nint   VSS     VSS     N   L=0.18U  W=0.83U  
M12     U35_out nint   VDD     VDD     P   L=0.18U  W=1.83U  
M13     u7_S    U35_out VSS     VSS     N   L=0.18U  W=0.83U  
M14     u7_S    U35_out VDD     VDD     P   L=0.184U  W=1.82U  
M15     SO      u3_in   VSS     VSS     N   L=0.18U  W=1.38U  
M16     SO      u3_in   VDD     VDD     P   L=0.184U  W=4.1U  
M17     u3_in   u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M18     u3_in   u9_D    VDD     VDD     P   L=0.18U  W=1.88U  
M19     u9_S    u3_in   VSS     VSS     N   L=0.18U  W=0.83U  
M20     u9_S    u3_in   VDD     VDD     P   L=0.185U  W=1.88U  
M21     U48_drain D       U48_source VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M22     U48_drain SD      U50_source VSS     N   L=0.18U  W=0.66U   
+  PS=.480U PD=.480U
M23     U50_source U71_out VSS     VSS     N   L=0.18U  W=0.66U
M24     U48_source U72_out VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M25     U81_drain U1_out  VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=1.164U
M26     U78_drain OE      U81_drain VSS     N   L=0.18U  W=0.69U   
+  PS=1.164U PD=1.239U
M27     U81_drain U35_out   VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=1.164U
M28     Z       U81_drain VSS     VSS     N   L=0.18U  W=1.38U   
+  PD=1.330U
M29     U66_drain SD      U48_drain VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M30     U67_drain D       U48_drain VDD     P   L=0.185U  W=1.78U   
+  PS=.520U PD=.520U
M31     VDD     U71_out U67_drain VDD     P   L=0.185U  W=1.78U   
+  PS=.520U
M32     VDD     U72_out U66_drain VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M33     U78_drain OE      VDD     VDD     P   L=0.184U  W=2.05U   
+  PD=1.227U
M34     Z       U78_drain VDD     VDD     P   L=0.182U  W=4.1U   
+  PD=2.018U
M35     U81_drain U1_out  U78_drain VDD     P   L=0.184U  W=2.05U   
+  PS=1.227U PD=1.145U
M36     U78_drain U35_out   VDD     VDD     P   L=0.18U  W=2.05U   
+  PD=1.227U
M37     U48_drain u10_out nint   VDD     P   L=0.18U  W=1.38U   
+  PD=.520U
M38     U48_drain u11_out nint   VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M39     u7_S    u11_out nint   VDD     P   L=0.18U  W=1.38U  
M40     u7_S    u10_out nint   VSS     N   L=0.18U  W=0.46U  
M41     u9_S    u10_out u9_D    VDD     P   L=0.18U  W=0.69U  
M42     u9_S    u11_out u9_D    VSS     N   L=0.18U  W=0.42U  
M43     U35_out u11_out u9_D    VDD     P   L=0.18U  W=0.69U  
M44     U35_out u10_out u9_D    VSS     N   L=0.18U  W=0.46U  

.ENDS slnht2

.SUBCKT slnht4 SO Z  D E OE SC SD VDD VSS
M1      U1_out  OE      VSS     VSS     N   L=0.18U  W=0.69U
M2      U1_out  OE      VDD     VDD     P   L=0.184U  W=2.05U
M3      U72_out SC      VSS     VSS     N   L=0.18U  W=0.69U
M4      U72_out SC      VDD     VDD     P   L=0.184U  W=1.91U
M5      U71_out U72_out VSS     VSS     N   L=0.18U  W=0.69U
M6      U71_out U72_out VDD     VDD     P   L=0.184U  W=1.91U
M7      u10_out E       VSS     VSS     N   L=0.18U  W=0.66U
M8      u10_out E       VDD     VDD     P   L=0.184U  W=1.74U
M9      u11_out u10_out VSS     VSS     N   L=0.18U  W=0.66U
M10     u11_out u10_out VDD     VDD     P   L=0.184U  W=1.74U
M11     U35_out nint   VSS     VSS     N   L=0.18U  W=0.83U
M12     U35_out nint   VDD     VDD     P   L=0.18U  W=1.83U
M13     u7_S    U35_out VSS     VSS     N   L=0.18U  W=0.83U
M14     u7_S    U35_out VDD     VDD     P   L=0.184U  W=1.83U
M15     SO      u3_in   VSS     VSS     N   L=0.18U  W=2.77U
M16     SO      u3_in   VDD     VDD     P   L=0.183U  W=8.20U
M17     u3_in   u9_D    VSS     VSS     N   L=0.18U  W=0.83U
M18     u3_in   u9_D    VDD     VDD     P   L=0.18U  W=1.88U
M19     u9_S    u3_in   VSS     VSS     N   L=0.18U  W=0.83U
M20     u9_S    u3_in   VDD     VDD     P   L=0.185U  W=1.88U
M21     U48_drain D       U48_source VSS     N   L=0.18U  W=0.69U
+  PS=.480U PD=.480U
M22     U48_drain SD      U50_source VSS     N   L=0.18U  W=0.66U
+  PS=.480U PD=.480U
M23     U50_source U71_out VSS     VSS     N   L=0.18U  W=0.66U
+  PD=.480U
M24     U48_source U72_out VSS     VSS     N   L=0.18U W=0.69U
+  PD=.480U
M25     U81_drain U1_out  VSS     VSS     N   L=0.18U  W=0.69U
+  PD=1.164U
M26     U78_drain OE      U81_drain VSS     N   L=0.18U  W=0.69U
+  PS=1.164U PD=1.239U
M27     U81_drain U35_out   VSS     VSS     N   L=0.18U  W=0.69U
+  PD=1.164U
M28     Z       U81_drain VSS     VSS     N   L=0.18U  W=2.77U
+  PD=1.330U
M29     U66_drain SD      U48_drain VDD     P   L=0.184U  W=1.91U
+  PS=.520U PD=.520U
M30     U67_drain D       U48_drain VDD     P   L=0.185U  W=1.78U
+  PS=.520U PD=.520U
M31     VDD     U71_out U67_drain VDD     P   L=0.185U  W=1.78U
+  PS=.520U
M32     VDD     U72_out U66_drain VDD     P   L=0.184U  W=1.91U
+  PS=.520U
M33     U78_drain OE      VDD     VDD     P   L=0.184U  W=2.05U
+  PD=1.227U
M34     Z       U78_drain VDD     VDD     P   L=0.182U  W=8.2U
+  PD=2.018U
M35     U81_drain U1_out  U78_drain VDD     P   L=0.184U  W=2.05U
+  PS=1.227U PD=1.145U
M36     U78_drain U35_out   VDD     VDD     P   L=0.18U  W=2.05U
+  PD=1.227U
M37     U48_drain u10_out nint   VDD     P   L=0.18U  W=1.38U
+  PD=.520U
M38     U48_drain u11_out nint   VSS     N   L=0.18U  W=0.46U
+  PD=.480U
M39     u7_S    u11_out nint   VDD     P   L=0.18U  W=1.38U
M40     u7_S    u10_out nint   VSS     N   L=0.18U  W=0.46U
M41     u9_S    u10_out u9_D    VDD     P   L=0.18U  W=0.73U
M42     u9_S    u11_out u9_D    VSS     N   L=0.18U  W=0.42U
M43     U35_out u11_out u9_D    VDD     P   L=0.18U  W=0.73U
M44     U35_out u10_out u9_D    VSS     N   L=0.18U  W=0.46U

.ENDS slnht4

.SUBCKT slnlb1 SO Q QN  D EN SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U      W=0.83U
M2      U35_out U35_in  VDD     VDD     P   L=0.185U     W=1.83U
M3      U37_out U35_out VSS     VSS     N   L=0.18U      W=0.83U
M4      U37_out U35_out VDD     VDD     P   L=0.186U      W=1.87U
M5      U38_out U38_in  VSS     VSS     N   L=0.18U      W=0.83U
M6      U38_out U38_in  VDD     VDD     P   L=0.184U      W=1.88U
M7      SO      U38_out VSS     VSS     N   L=0.18U      W=0.69U
M8      SO      U38_out VDD     VDD     P   L=0.184U      W=2.05U
M9      U15_G   EN      VSS     VSS     N   L=0.18U      W=0.66U
M10     U15_G   EN      VDD     VDD     P   L=0.184U      W=1.74U
M11     U15_GB  U15_G   VSS     VSS     N   L=0.18U      W=0.66U
M12     U15_GB  U15_G   VDD     VDD     P   L=0.184U      W=1.74U
M13     U43_gate U45_gate VSS     VSS     N   L=0.18U     W=0.69U
M14     U43_gate U45_gate VDD     VDD     P   L=0.184U      W=1.91U
M15     U45_gate SC      VSS     VSS     N   L=0.18U      W=0.69U
M16     U45_gate SC      VDD     VDD     P   L=0.184U      W=1.91U
M17     u9_S    U38_out VSS     VSS     N   L=0.18U      W=0.83U
M18     u9_S    U38_out VDD     VDD     P   L=0.184U      W=1.88U
M19     QN      U35_out VSS     VSS     N   L=0.18U      W=0.69U
M20     QN      U35_out VDD     VDD     P   L=0.184U      W=2.05U
M21     Q       U35_in  VSS     VSS     N   L=0.18U      W=0.69U
M22     Q       U35_in  VDD     VDD     P   L=0.184U      W=2.05U
M23     U66_drain SD      U66_source VDD     P   L=0.184U       W=1.91U
+  PS=.520U PD=.520U
M24     VDD     U45_gate U66_drain VDD     P   L=0.184U       W=1.91U
+  PS=.520U
M25     VDD     U43_gate U43_source VDD     P   L=0.184U       W=1.78U
+  PS=.520U
M26     U43_source D       U66_source VDD     P   L=0.184U       W=1.78U
+  PS=.520U PD=.520U
M27     U66_source U15_GB  U35_in  VDD     P   L=0.185U       W=1.44U
+  PD=.520U
M28     U66_source U15_G   U35_in  VSS     N   L=0.18U       W=0.46U
+  PD=.480U
M29     U35_out U15_G   U38_in  VDD     P   L=0.18U      W=0.69U
M30     U35_out U15_GB  U38_in  VSS     N   L=0.18U      W=0.46U
M31     U37_out U15_G   U35_in  VDD     P   L=0.18U      W=1.44U
M32     U37_out U15_GB  U35_in  VSS     N   L=0.18U      W=0.46U
M33     u9_S    U15_GB  U38_in  VDD     P   L=0.18U      W=0.69U
M34     u9_S    U15_G   U38_in  VSS     N   L=0.18U      W=0.42U
M35     U68_drain U45_gate VSS     VSS     N   L=0.18U       W=0.69U
+  PD=.480U
M36     U66_source D       U68_drain VSS     N   L=0.18U       W=0.69U
+  PS=.480U PD=.480U
M37     U69_drain U43_gate VSS     VSS     N   L=0.18U       W=0.66U
+  PD=.480U
M38     U66_source SD      U69_drain VSS     N   L=0.18U       W=0.66U
+  PS=.480U PD=.480U

.ENDS slnlb1

.SUBCKT slnlb2 SO Q QN  D EN SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U      W=0.83U
M2      U35_out U35_in  VDD     VDD     P   L=0.184U      W=1.83U
M3      U37_out U35_out VSS     VSS     N   L=0.18U      W=0.83U
M4      U37_out U35_out VDD     VDD     P   L=0.185U     W=1.83U
M5      U38_out U38_in  VSS     VSS     N   L=0.18U     W=0.83U
M6      U38_out U38_in  VDD     VDD     P   L=0.184U      W=1.88U
M7      SO      U38_out VSS     VSS     N   L=0.18U     W=1.38U
M8      SO      U38_out VDD     VDD     P   L=0.182U      W=4.10U
M9      U15_G   EN      VSS     VSS     N   L=0.18U      W=0.66U
M10     U15_G   EN      VDD     VDD     P   L=0.184U      W=1.74U
M11     U15_GB  U15_G   VSS     VSS     N   L=0.18U     W=0.66U
M12     U15_GB  U15_G   VDD     VDD     P   L=0.184U     W=1.74U
M13     U43_gate U45_gate VSS     VSS     N   L=0.18U      W=0.69U
M14     U43_gate U45_gate VDD     VDD     P   L=0.184U     W=1.91U
M15     U45_gate SC      VSS     VSS     N   L=0.18U      W=0.69U
M16     U45_gate SC      VDD     VDD     P   L=0.184U     W=1.91U
M17     u9_S    U38_out VSS     VSS     N   L=0.18U      W=0.83U
M18     u9_S    U38_out VDD     VDD     P   L=0.184U      W=1.88U
M19     QN      U35_out VSS     VSS     N   L=0.185U     W=1.38U
M20     QN      U35_out VDD     VDD     P   L=0.182U     W=4.10U
M21     Q       U35_in  VSS     VSS     N   L=0.185U      W=1.38U
M22     Q       U35_in  VDD     VDD     P   L=0.184U      W=4.10U
M23     U66_drain SD      U66_source VDD     P   L=0.184U      W=1.91U
+  PS=.520U PD=.520U
M24     VDD     U45_gate U66_drain VDD     P   L=0.184U       W=1.91U
+  PS=.520U
M25     VDD     U43_gate U43_source VDD     P   L=0.184U       W=1.78U
+  PS=.520U
M26     U43_source D       U66_source VDD     P   L=0.184U       W=1.78U
+  PS=.520U PD=.520U
M27     U66_source U15_GB  U35_in  VDD     P   L=0.185U       W=1.44U
+  PD=.520U
M28     U66_source U15_G   U35_in  VSS     N   L=0.18U       W=0.46U
+  PD=.480U
M29     U35_out U15_G   U38_in  VDD     P   L=0.18U      W=0.69U
M30     U35_out U15_GB  U38_in  VSS     N   L=0.18U      W=0.46U
M31     U37_out U15_G   U35_in  VDD     P   L=0.18U      W=1.44U
M32     U37_out U15_GB  U35_in  VSS     N   L=0.18U      W=0.46U
M33     u9_S    U15_GB  U38_in  VDD     P   L=0.18U     W=0.69U
M34     u9_S    U15_G   U38_in  VSS     N   L=0.18U      W=0.42U
M35     U68_drain U45_gate VSS     VSS     N   L=0.18U       W=0.69U
+  PD=.480U
M36     U66_source D       U68_drain VSS     N   L=0.18U       W=0.69U
+  PS=.480U PD=.480U
M37     U69_drain U43_gate VSS     VSS     N   L=0.18U       W=0.66U
+  PD=.480U
M38     U66_source SD      U69_drain VSS     N   L=0.18U       W=0.66U
+  PS=.480U PD=.480U

.ENDS slnlb2

.SUBCKT slnlb4 SO Q QN  D EN SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U     W=0.83U
M2      U35_out U35_in  VDD     VDD     P   L=0.184U      W=1.83U
M3      U37_out U35_out VSS     VSS     N   L=0.18U      W=0.83U
M4      U37_out U35_out VDD     VDD     P   L=0.185U     W=1.83U
M5      U38_out U38_in  VSS     VSS     N   L=0.18U      W=0.83U
M6      U38_out U38_in  VDD     VDD     P   L=0.184U      W=1.88U
M7      SO      U38_out VSS     VSS     N   L=0.18U      W=2.77U
M8      SO      U38_out VDD     VDD     P   L=0.182U      W=8.20U
M9      U15_G   EN      VSS     VSS     N   L=0.18U      W=0.66U
M10     U15_G   EN      VDD     VDD     P   L=0.184U      W=1.74U
M11     U15_GB  U15_G   VSS     VSS     N   L=0.18U      W=0.66U
M12     U15_GB  U15_G   VDD     VDD     P   L=0.184U      W=1.74U
M13     U43_gate U45_gate VSS     VSS     N   L=0.18U      W=0.69U
M14     U43_gate U45_gate VDD     VDD     P   L=0.184U      W=1.91U
M15     U45_gate SC      VSS     VSS     N   L=0.18U      W=0.69U
M16     U45_gate SC      VDD     VDD     P   L=0.184U     W=1.91U
M17     u9_S    U38_out VSS     VSS     N   L=0.18U      W=0.83U
M18     u9_S    U38_out VDD     VDD     P   L=0.184U      W=1.88U
M19     QN      U35_out VSS     VSS     N   L=0.18U      W=2.77U
M20     QN      U35_out VDD     VDD     P   L=0.182U      W=8.20U
M21     Q       U35_in  VSS     VSS     N   L=0.18U     W=2.77U
M22     Q       U35_in  VDD     VDD     P   L=0.18U     W=8.20U
M23     U66_drain SD      U66_source VDD     P   L=0.184U       W=1.91U
+  PS=.520U PD=.520U
M24     VDD     U45_gate U66_drain VDD     P   L=0.184U       W=1.91U
+  PS=.520U
M25     VDD     U43_gate U43_source VDD     P   L=0.184U       W=1.78U
+  PS=.520U
M26     U43_source D       U66_source VDD     P   L=0.184U       W=1.78U
+  PS=.520U PD=.520U
M27     U66_source U15_GB  U35_in  VDD     P   L=0.185U       W=1.44U
+  PD=.520U
M28     U66_source U15_G   U35_in  VSS     N   L=0.18U      W=0.46U
+  PD=.480U
M29     U35_out U15_G   U38_in  VDD     P   L=0.18U      W=0.69U
M30     U35_out U15_GB  U38_in  VSS     N   L=0.18U      W=0.46U
M31     U37_out U15_G   U35_in  VDD     P   L=0.18U      W=1.44U
M32     U37_out U15_GB  U35_in  VSS     N   L=0.18U      W=0.46U
M33     u9_S    U15_GB  U38_in  VDD     P   L=0.18U     W=0.69U
M34     u9_S    U15_G   U38_in  VSS     N   L=0.18U      W=0.42U
M35     U68_drain U45_gate VSS     VSS     N   L=0.18U    W=0.69U
+  PD=.480U
M36     U66_source D       U68_drain VSS     N   L=0.18U      W=0.69U
+  PS=.480U PD=.480U
M37     U69_drain U43_gate VSS     VSS     N   L=0.18U      W=0.66U
+  PD=.480U
M38     U66_source SD      U69_drain VSS     N   L=0.18U     W=0.66U
+  PS=.480U PD=.480U

.ENDS slnlb4

.SUBCKT slnln1 SO QN  D EN SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.83U  
M2      U35_out U35_in  VDD     VDD     P   L=0.185U  W=1.83U  
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.83U  
M4      U37_out U35_out VDD     VDD     P   L=0.18U  W=1.83U  
M5      u7_GB   EN      VSS     VSS     N   L=0.18U  W=0.66U  
M6      u7_GB   EN      VDD     VDD     P   L=0.18U  W=1.74U  
M7      u7_G    u7_GB   VSS     VSS     N   L=0.18U  W=0.66U  
M8      u7_G    u7_GB   VDD     VDD     P   L=0.18U  W=1.74U  
M9      U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U  
M10     U43_gate U68_gate VDD     VDD     P   L=0.18U  W=1.91U  
M11     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M12     U68_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M13     u9_S    U36_in  VSS     VSS     N   L=0.18U  W=.83U  
M14     u9_S    U36_in  VDD     VDD     P   L=0.184U  W=1.88U  
M15     U36_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M16     U36_in  u9_D    VDD     VDD     P   L=0.185U  W=1.88U  
M17     SO      U36_in  VSS     VSS     N   L=0.18U  W=0.69U  
M18     SO      U36_in  VDD     VDD     P   L=0.186U  W=1.95U  
M19     QN      U35_out VSS     VSS     N   L=0.18U  W=0.69U  
M20     QN      U35_out VDD     VDD     P   L=0.186U  W=1.94U  
M21     VDD     U43_gate U43_source VDD     P   L=0.18U  W=1.78U   
+  PS=.520U
M22     U43_source D       U67_source VDD     P   L=0.18U  W=1.78U   
+  PS=.520U PD=.520U
M23     VDD     U68_gate U45_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M24     U45_source SD      U67_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M25     U68_drain U68_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M26     U67_source D       U68_drain VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M27     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M28     U67_source SD      U69_drain VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U
M29     U37_out u7_GB   U35_in  VDD     P   L=0.185U  W=1.44U  
M30     U37_out u7_G    U35_in  VSS     N   L=0.18U  W=0.46U  
M31     U67_source u7_G    U35_in  VDD     P   L=0.18U  W=1.44U   
+  PD=.520U
M32     U67_source u7_GB   U35_in  VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M33     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.69U  
M34     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M35     U35_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.69U  
M36     U35_out u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  

.ENDS slnln1

.SUBCKT slnln2 SO QN  D EN SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.83U
M2      U35_out U35_in  VDD     VDD     P   L=0.18U  W=1.83U
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.83U
M4      U37_out U35_out VDD     VDD     P   L=0.184U  W=1.83U
M5      u7_GB   EN      VSS     VSS     N   L=0.18U  W=0.66U
M6      u7_GB   EN      VDD     VDD     P   L=0.184U  W=1.74U
M7      u7_G    u7_GB   VSS     VSS     N   L=0.18U  W=0.66U
M8      u7_G    u7_GB   VDD     VDD     P   L=0.184U  W=1.74U
M9      U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U
M10     U43_gate U68_gate VDD     VDD     P   L=0.18U  W=1.91U
M11     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U
M12     U68_gate SC      VDD     VDD     P   L=0.184U  W=1.91U
M13     u9_S    U36_in  VSS     VSS     N   L=0.18U  W=0.83U
M14     u9_S    U36_in  VDD     VDD     P   L=0.18U  W=1.88U
M15     U36_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U
M16     U36_in  u9_D    VDD     VDD     P   L=0.185U  W=1.88U
M17     SO      U36_in  VSS     VSS     N   L=0.18U  W=1.38U
M18     SO      U36_in  VDD     VDD     P   L=0.183U  W=4.10U
M19     QN      U35_out VSS     VSS     N   L=0.18U  W=1.38U
M20     QN      U35_out VDD     VDD     P   L=0.18U  W=4.10U
M21     VDD     U43_gate U43_source VDD     P   L=0.18U  W=1.78U
+  PS=.520U
M22     U43_source D       U67_source VDD     P   L=0.18U  W=1.78U
+  PS=.520U PD=.520U
M23     VDD     U68_gate U45_source VDD     P   L=0.184U  W=1.91U
+  PS=.520U
M24     U45_source SD      U67_source VDD     P   L=0.184U  W=1.91U
+  PS=.520U PD=.520U
M25     U68_drain U68_gate VSS     VSS     N   L=0.18U  W=0.69U
+  PD=.480U
M26     U67_source D       U68_drain VSS     N   L=0.18U  W=0.69U
+  PS=.480U PD=.480U
M27     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=0.66U
+  PD=.480U
M28     U67_source SD      U69_drain VSS     N   L=0.18U  W=0.66U
+  PS=.480U PD=.480U
M29     U37_out u7_GB   U35_in  VDD     P   L=0.18U  W=1.44U
M30     U37_out u7_G    U35_in  VSS     N   L=0.18U  W=0.46U
M31     U67_source u7_G    U35_in  VDD     P   L=0.18U  W=1.44U
+  PD=.520U
M32     U67_source u7_GB   U35_in  VSS     N   L=0.18U  W=0.46U
+  PD=.480U
M33     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.69U
M34     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U
M35     U35_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.69U
M36     U35_out u7_G    u9_D    VSS     N   L=0.18U  W=0.46U

.ENDS slnln2

.SUBCKT slnln4 SO QN  D EN SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS     N   L=0.18U  W=0.83U  
M2      U35_out U35_in  VDD     VDD     P   L=0.185U  W=1.83U  
M3      U37_out U35_out VSS     VSS     N   L=0.18U  W=0.83U  
M4      U37_out U35_out VDD     VDD     P   L=0.18U  W=1.83U  
M5      u7_GB   EN      VSS     VSS     N   L=0.18U  W=0.66U  
M6      u7_GB   EN      VDD     VDD     P   L=0.18U  W=1.74U  
M7      u7_G    u7_GB   VSS     VSS     N   L=0.18U  W=0.66U  
M8      u7_G    u7_GB   VDD     VDD     P   L=0.18U  W=1.74U  
M9      U43_gate U68_gate VSS     VSS     N   L=0.18U  W=0.69U  
M10     U43_gate U68_gate VDD     VDD     P   L=0.18U  W=1.91U  
M11     U68_gate SC      VSS     VSS     N   L=0.18U  W=0.69U  
M12     U68_gate SC      VDD     VDD     P   L=0.184U  W=1.91U  
M13     u9_S    U36_in  VSS     VSS     N   L=0.18U  W=.83U  
M14     u9_S    U36_in  VDD     VDD     P   L=0.184U  W=1.88U  
M15     U36_in  u9_D    VSS     VSS     N   L=0.18U  W=0.83U  
M16     U36_in  u9_D    VDD     VDD     P   L=0.185U  W=1.88U  
M17     SO      U36_in  VSS     VSS     N   L=0.18U  W=2.77U  
M18     SO      U36_in  VDD     VDD     P   L=0.187U  W=8.2U  
M19     QN      U35_out VSS     VSS     N   L=0.18U  W=2.77U  
M20     QN      U35_out VDD     VDD     P   L=0.184U  W=8.2U  
M21     VDD     U43_gate U43_source VDD     P   L=0.18U  W=1.78U   
+  PS=.520U
M22     U43_source D       U67_source VDD     P   L=0.18U  W=1.78U   
+  PS=.520U PD=.520U
M23     VDD     U68_gate U45_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U
M24     U45_source SD      U67_source VDD     P   L=0.184U  W=1.91U   
+  PS=.520U PD=.520U
M25     U68_drain U68_gate VSS     VSS     N   L=0.18U  W=0.69U   
+  PD=.480U
M26     U67_source D       U68_drain VSS     N   L=0.18U  W=0.69U   
+  PS=.480U PD=.480U
M27     U69_drain U43_gate VSS     VSS     N   L=0.18U  W=.66U   
+  PD=.480U
M28     U67_source SD      U69_drain VSS     N   L=0.18U  W=.66U   
+  PS=.480U PD=.480U
M29     U37_out u7_GB   U35_in  VDD     P   L=0.185U  W=1.44U  
M30     U37_out u7_G    U35_in  VSS     N   L=0.18U  W=0.46U  
M31     U67_source u7_G    U35_in  VDD     P   L=0.18U  W=1.44U   
+  PD=.520U
M32     U67_source u7_GB   U35_in  VSS     N   L=0.18U  W=0.46U   
+  PD=.480U
M33     u9_S    u7_G    u9_D    VDD     P   L=0.18U  W=0.69U  
M34     u9_S    u7_GB   u9_D    VSS     N   L=0.18U  W=0.42U  
M35     U35_out u7_GB   u9_D    VDD     P   L=0.18U  W=0.69U  
M36     U35_out u7_G    u9_D    VSS     N   L=0.18U  W=0.46U  

.ENDS slnln4

.SUBCKT slnlq1 SO Q  D EN SC SD VDD VSS
M1      U35_out U35_in  VSS       VSS     N   L=0.18U       W=0.83U
M2      U35_out U35_in  VDD       VDD     P   L=0.18U       W=1.83U
M3      U37_out U35_out VSS       VSS     N   L=0.18U       W=0.83U
M4      U37_out U35_out VDD       VDD     P   L=0.18U       W=1.83U
M5      U38_out u8_D    VSS       VSS     N   L=0.18U       W=0.83U
M6      U38_out u8_D    VDD       VDD     P   L=0.18U       W=1.88U
M7      SO      U38_out VSS       VSS     N   L=0.18U       W=0.69U
M8      SO      U38_out VDD       VDD     P   L=0.184U      W=2.05U
M9      U15_G   EN      VSS         VSS     N   L=0.18U       W=0.66U
M10     U15_G   EN      VDD         VDD     P   L=0.184U      W=1.74U
M11     U15_GB  U15_G   VSS         VSS     N   L=0.18U       W=0.66U
M12     U15_GB  U15_G   VDD         VDD     P   L=0.18U       W=1.74U
M13     U43_gate U45_gate VSS       VSS     N   L=0.18U       W=0.69U
M14     U43_gate U45_gate VDD       VDD     P   L=0.18U       W=1.91U
M15     U45_gate SC      VSS        VSS     N   L=0.18U       W=0.69U
M16     U45_gate SC      VDD        VDD     P   L=0.184U      W=1.91U
M17     U36_out U38_out VSS         VSS     N   L=0.18U       W=0.83U
M18     U36_out U38_out VDD         VDD     P   L=0.184U      W=1.88U
M19     Q       U35_in  VSS         VSS     N   L=0.18U       W=0.69U
M20     Q       U35_in  VDD         VDD     P   L=0.187U      W=2.01U
M21     U15_S   U15_GB  U35_in      VDD     P   L=0.18U   PD=.520U    W=1.44U
M22     U15_S   U15_G   U35_in      VSS     N   L=0.18U   PD=.480U    W=0.46U
M23     U37_out U15_G   U35_in      VDD     P   L=0.186U      W=1.44U
M24     U37_out U15_GB  U35_in      VSS     N   L=0.18U       W=0.46U
M25     U35_out U15_G   u8_D        VDD     P   L=0.18U       W=0.69U
M26     U35_out U15_GB  u8_D        VSS     N   L=0.18U       W=0.46U
M27     U36_out U15_GB  u8_D        VDD     P   L=0.18U       W=0.69U
M28     U36_out U15_G   u8_D        VSS     N   L=0.18U       W=0.42U
M29     U66_drain SD      U15_S     VDD     P   L=0.18U       W=1.91U
+  PS=.520U PD=.520U
M30     VDD     U45_gate U66_drain  VDD     P   L=0.18U       W=1.91U
+  PS=.520U
M31     VDD     U43_gate U43_source VDD     P   L=0.185U      W=1.78U
+  PS=.520U
M32     U43_source D       U15_S    VDD     P   L=0.185U      W=1.78U
+  PS=.520U PD=.520U
M33     U68_drain U45_gate VSS      VSS     N   L=0.18U       W=0.69U
+  PD=.480U
M34     U15_S   D       U68_drain   VSS     N   L=0.18U       W=0.69U
+  PS=.480U PD=.480U
M35     U69_drain U43_gate VSS      VSS     N   L=0.18U       W=0.66U
+  PD=.480U
M36     U15_S   SD      U69_drain   VSS     N   L=0.18U       W=0.66U
+  PS=.480U PD=.480U

.ENDS slnlq1

.SUBCKT slnlq2 SO Q  D EN SC SD VDD VSS
M1      U35_out U35_in  VSS     VSS       N   L=0.18U      W=0.83U
M2      U35_out U35_in  VDD     VDD       P   L=0.18U      W=1.83U
M3      U37_out U35_out VSS     VSS       N   L=0.18U      W=0.83U
M4      U37_out U35_out VDD     VDD       P   L=0.185U     W=1.74U
M5      U38_out u8_D    VSS     VSS       N   L=0.18U      W=0.83U
M6      U38_out u8_D    VDD     VDD       P   L=0.18U      W=1.88U
M7      SO      U38_out VSS     VSS       N   L=0.186U     W=1.38U
M8      SO      U38_out VDD     VDD       P   L=0.184U     W=4.099U
M9      U15_G   EN      VSS     VSS       N   L=0.18U      W=0.66U
M10     U15_G   EN      VDD     VDD       P   L=0.184U     W=1.74U
M11     U15_GB  U15_G   VSS     VSS       N   L=0.18U      W=0.66U
M12     U15_GB  U15_G   VDD     VDD       P   L=0.18U      W=1.74U
M13     U43_gate U45_gate VSS     VSS     N   L=0.18U      W=0.69U
M14     U43_gate U45_gate VDD     VDD     P   L=0.18U      W=1.91U
M15     U45_gate SC      VSS     VSS      N   L=0.18U      W=0.69U
M16     U45_gate SC      VDD     VDD      P   L=0.184U     W=1.91U
M17     U36_out U38_out VSS     VSS       N   L=0.18U      W=0.83U
M18     U36_out U38_out VDD     VDD       P   L=0.184U     W=1.88U
M19     Q       U35_in  VSS     VSS       N   L=0.18U      W=1.38U
M20     Q       U35_in  VDD     VDD       P   L=0.186U     W=3.87U
M21     U15_S   U15_GB  U35_in  VDD       P   L=0.18U     PD=.520U  W=1.44U
M22     U15_S   U15_G   U35_in  VSS       N   L=0.18U     PD=.480U  W=0.46U
M23     U37_out U15_G   U35_in  VDD       P   L=0.186U     W=1.44U
M24     U37_out U15_GB  U35_in  VSS       N   L=0.18U      W=0.46U
M25     U35_out U15_G   u8_D    VDD       P   L=0.18U      W=0.69U
M26     U35_out U15_GB  u8_D    VSS       N   L=0.18U      W=0.46U
M27     U36_out U15_GB  u8_D    VDD       P   L=0.18U      W=0.69U
M28     U36_out U15_G   u8_D    VSS       N   L=0.18U      W=0.42U
M29     U66_drain SD      U15_S   VDD     P   L=0.18U      W=1.91U
+  PS=.520U PD=.520U
M30     VDD     U45_gate U66_drain VDD    P   L=0.18U      W=1.91U
+  PS=.520U
M31     VDD     U43_gate U43_source VDD   P   L=0.185U     W=1.78U
+  PS=.520U
M32     U43_source D       U15_S   VDD    P   L=0.185U     W=1.78U
+  PS=.520U PD=.520U
M33     U68_drain U45_gate VSS     VSS    N   L=0.18U      W=0.69U
+  PD=.480U
M34     U15_S   D       U68_drain VSS     N   L=0.18U      W=0.69U
+  PS=.480U PD=.480U
M35     U69_drain U43_gate VSS     VSS    N   L=0.18U      W=0.66U
+  PD=.480U
M36     U15_S   SD      U69_drain VSS     N   L=0.18U      W=0.66U
+  PS=.480U PD=.480U

.ENDS slnlq2

.SUBCKT slnlq4 SO Q  D EN SC SD VDD VSS
M1      U35_out U35_in  VSS       VSS         N   L=0.18U        W=0.83U
M2      U35_out U35_in  VDD       VDD         P   L=0.18U        W=1.83U
M3      U37_out U35_out VSS       VSS         N   L=0.18U        W=0.83U
M4      U37_out U35_out VDD       VDD         P   L=0.185U       W=1.83U
M5      U38_out U38_in  VSS       VSS         N   L=0.18U        W=0.83U
M6      U38_out U38_in  VDD       VDD         P   L=0.184U       W=1.88U
M7      SO      U38_out VSS       VSS         N   L=0.183U       W=2.77U
M8      SO      U38_out VDD       VDD         P   L=0.184U       W=8.197U
M9      u8_GB   EN      VSS       VSS         N   L=0.18U        W=0.66U
M10     u8_GB   EN      VDD       VDD         P   L=0.185U       W=1.74U
M11     u8_G    u8_GB   VSS       VSS         N   L=0.18U        W=0.66U
M12     u8_G    u8_GB   VDD       VDD         P   L=0.18U        W=1.74U
M13     U43_gate U45_gate VSS     VSS         N   L=0.18U        W=0.69U
M14     U43_gate U45_gate VDD     VDD         P   L=0.18U        W=1.91U
M15     U45_gate SC      VSS      VSS         N   L=0.18U        W=0.69U
M16     U45_gate SC      VDD      VDD         P   L=0.184U       W=1.91U
M17     u9_S    U38_out VSS       VSS         N   L=0.18U        W=0.83U
M18     u9_S    U38_out VDD       VDD         P   L=0.184U       W=1.88U
M19     Q       U35_in  VSS       VSS         N   L=0.18U        W=2.77U
M20     Q       U35_in  VDD       VDD         P   L=0.18975U     W=8.1969U
M21     U66_drain SD      U66_source VDD      P   L=0.18U        W=1.91U
+  PS=.520U PD=.520U
M22     VDD     U45_gate U66_drain VDD        P   L=0.18U        W=1.91U
+  PS=.520U
M23     VDD     U43_gate U43_source VDD       P   L=0.185U       W=1.78U
+  PS=.520U
M24     U43_source D       U66_source VDD     P   L=0.185U       W=1.78U
+  PS=.520U PD=.520U
M25     U68_drain U45_gate VSS     VSS        N   L=0.18U        W=0.69U
+  PD=.480U
M26     U66_source D       U68_drain VSS      N   L=0.18U        W=0.69U
+  PS=.480U PD=.480U
M27     U69_drain U43_gate VSS     VSS        N   L=0.18U        W=0.66U
+  PD=.480U
M28     U66_source SD      U69_drain VSS      N   L=0.18U        W=0.66U
+  PS=.480U PD=.480U
M29     U35_out u8_GB   U38_in  VDD           P   L=0.18U        W=0.69U
M30     U35_out u8_G    U38_in  VSS           N   L=0.18U        W=0.46U
M31     U37_out u8_GB   U35_in  VDD           P   L=0.186U       W=1.44U
M32     U37_out u8_G    U35_in  VSS           N   L=0.18U        W=0.46U
M33     U66_source u8_G    U35_in  VDD        P   L=0.18U        W=1.44U
+  PD=.520U
M34     U66_source u8_GB   U35_in  VSS        N   L=0.18U        W=0.46U
+  PD=.480U
M35     u9_S    u8_G    U38_in  VDD           P   L=0.18U        W=0.69U
M36     u9_S    u8_GB   U38_in  VSS           N   L=0.18U        W=0.42U

.ENDS slnlq4

.SUBCKT srlab4 Q QN  RN SN VDD VSS
M1      U6_u7_drain SN      VSS     VSS     N   L=0.18U      W=0.92U
M2      U6_out  U6_in1  U6_u7_drain VSS     N   L=0.18U      W=0.92U
M3      U6_out  U6_in1  VDD     VDD     P   L=0.185U          W=1.66U
M4      VDD     SN      U6_out  VDD     P   L=0.18U          W=1.66U
M5      U7_u7_drain U6_out  VSS     VSS     N   L=0.18U      W=0.92U
M6      U6_in1  RN      U7_u7_drain VSS     N   L=0.18U      W=0.92U
M7      U6_in1  RN      VDD     VDD     P   L=0.185U          W=1.66U
M8      VDD     U6_out  U6_in1  VDD     P   L=0.18U          W=1.66U
M9      Q       U6_in1  VSS     VSS     N   L=0.18U          W=2.91U
M10     Q       U6_in1  VDD     VDD     P   L=0.184U          W=8.2U
M11     QN      U6_out  VSS     VSS     N   L=0.186U          W=2.91U
M12     QN      U6_out  VDD     VDD     P   L=0.184U          W=8.2U

.ENDS srlab4

.SUBCKT su01d4 CO S  A B CI VDD VSS
M1      U42_drain A       U42_source VDD     P   L=0.18U  W=1.34U
M2      U36_drain U36_gate VDD     VDD     P   L=0.18U  W=1.43U
M3      U38_drain CI      U38_source VDD     P   L=0.185U  W=1.43U
M4      U42_source U36_gate VDD     VDD     P   L=0.18U  W=1.34U
M5      U35_drain U36_gate VDD     VDD     P   L=0.185U  W=1.52U
M6      U38_source A       U36_drain VDD     P   L=0.185U  W=1.43U
M7      U42_drain CI      U32_source VDD     P   L=0.185U  W=1.56U
M8      U32_source U36_gate VDD     VDD     P   L=0.18U      W=1.56U
M9      U32_source A       VDD     VDD     P   L=0.185U      W=1.56U
M10     U35_drain CI      VDD     VDD     P   L=0.185U      W=1.52U
M11     U38_drain U42_drain U35_drain VDD     P   L=0.185U      W=1.43U
M12     U35_drain A       VDD     VDD     P   L=0.18U      W=1.56U
M13     U56_drain U36_gate VSS     VSS     N   L=0.18U      W=0.61U
M14     U48_drain U36_gate VSS     VSS     N   L=0.18U      W=0.61U
M15     U52_drain U36_gate VSS     VSS     N   L=0.18U      W=0.55U
M16     U51_drain A       U52_drain VSS     N   L=0.18U      W=0.55U
M17     U42_drain A       U48_drain VSS     N   L=0.18U      W=0.61U
M18     U47_drain U36_gate VSS     VSS     N   L=0.18U      W=0.61U
M19     U42_drain CI      U47_drain VSS     N   L=0.18U      W=0.61U
M20     U47_drain A       VSS     VSS     N   L=0.18U      W=0.61U
M21     U56_drain CI      VSS     VSS     N   L=0.18U      W=0.55U
M22     U38_drain U42_drain U56_drain VSS     N   L=0.18U      W=0.55U
M23     U56_drain A       VSS     VSS     N   L=0.18U      W=0.61U
M24     U38_drain CI      U51_drain VSS     N   L=0.18U      W=0.55U
M25     U36_gate B       VSS     VSS     N   L=0.18U      W=0.46U
M26     U36_gate B       VDD     VDD     P   L=0.186U      W=1.32U
M27     CO      U42_drain VSS     VSS     N   L=0.182U      W=2.91U
M28     CO      U42_drain VDD     VDD     P   L=0.182U      W=8.20U
M29     S       U38_drain VSS     VSS     N   L=0.182U      W=2.91U
M30     S       U38_drain VDD     VDD     P   L=0.182U      W=7.89U

.ENDS su01d4

.SUBCKT xn02d7 ZN  A1 A2 VDD VSS
M1      U7_drain   A2          VDD       VDD     P   L=0.18U   W=1.95U   
+  PD=1.589U
M2      U8_drain   A1          U7_drain  VDD     P   L=0.18U   W=1.95U   
+  PS=1.589U PD=1.555U
M3      U4_drain   U10_gate    VDD       VDD     P   L=0.183U  W=1.95U   
+  PD=1.520U
M4      U8_drain   U112_out    U4_drain  VDD     P   L=0.183U  W=1.95U   
+  PS=1.520U PD=1.555U
M5      U10_drain  U10_gate    VSS       VSS     N   L=0.18U   W=0.71U   
+  PD=1.025U
M6      U8_drain   A1          U10_drain VSS     N   L=0.18U   W=0.71U   
+  PS=1.025U PD=1.275U
M7      U8_drain   U112_out    U5_source VSS     N   L=0.18U   W=0.71U   
+  PS=1.524U PD=1.275U 
M8      U5_source  A2          VSS       VSS     N   L=0.18U   W=0.71U   
+  PD=1.524U
M9      ZN         U113_in     VSS       VSS     N   L=0.186U  W=5.05U  
M10     ZN         U113_in     VDD       VDD     P   L=0.182U  W=14.34U  
M11     U113_in    U8_drain    VSS       VSS     N   L=0.18U   W=1.69U  
M12     U113_in    U8_drain    VDD       VDD     P   L=0.184U  W=4.51U  
M13     U112_out   A1          VSS       VSS     N   L=0.18U   W=0.42U  
M14     U112_out   A1          VDD       VDD     P   L=0.186U  W=1.19U  
M15     U10_gate   A2          VSS       VSS     N   L=0.18U   W=0.42U  
M16     U10_gate   A2          VDD       VDD     P   L=0.186U  W=1.19U  

.ENDS xn02d7

.SUBCKT xn02da ZN  A1 A2 VDD VSS
M1      U7_drain  A2        VDD        VDD     P   L=0.18U   W=1.95U   
+  PD=1.589U 
M2      U8_drain  A1        U7_drain   VDD     P   L=0.18U   W=1.95U   
+  PS=1.589U PD=1.555U
M3      U4_drain  U10_gate  VDD        VDD     P   L=0.183U  W=1.95U   
+  PD=1.520U
M4      U8_drain  U112_out  U4_drain   VDD     P   L=0.183U  W=1.95U   
+  PS=1.520U PD=1.555U
M5      U10_drain U10_gate  VSS        VSS     N   L=0.18U   W=0.71U   
+  PD=1.025U
M6      U8_drain  A1        U10_drain  VSS     N   L=0.18U   W=0.71U   
+  PS=1.025U PD=1.275U 
M7      U8_drain  U112_out  U5_source  VSS     N   L=0.18U   W=0.71U   
+  PS=1.524U PD=1.275U
M8      U5_source A2        VSS        VSS     N   L=0.18U   W=0.71U   
+  PD=1.524U
M9      ZN        U113_in   VSS        VSS     N   L=0.187U  W=7.17U  
M10     ZN        U113_in   VDD        VDD     P   L=0.183U  W=20.49U  
M11     U113_in   U8_drain  VSS        VSS     N   L=0.183U  W=1.61U  
M12     U113_in   U8_drain  VDD        VDD     P   L=0.184U  W=4.51U  
M13     U112_out  A1        VSS        VSS     N   L=0.18U   W=0.42U  
M14     U112_out  A1        VDD        VDD     P   L=0.186U  W=1.19U  
M15     U10_gate  A2        VSS        VSS     N   L=0.18U   W=0.42U  
M16     U10_gate  A2        VDD        VDD     P   L=0.186U  W=1.19U  

.ENDS xn02da

.SUBCKT xr02d7 Z  A1 A2 VDD VSS
M1      U9_drain U9_gate U9_source VSS     N   L=0.18U  W=0.54U   
+  PS=.745U PD=.697U
M2      U9_source U10_gate VSS     VSS     N   L=0.18U  W=0.54U   
+  PD=.745U
M3      U63_drain A2      VSS     VSS     N   L=0.18U  W=0.54U   
+  PD=.613U
M4      U9_drain A1      U63_drain VSS     N   L=0.18U  W=0.54U   
+  PS=.613U PD=.697U
M5      Z       U195_gate VSS     VSS     N   L=0.18U  W=5.05U   
+  PD=1.069U
M6      U195_gate U9_drain VSS     VSS     N   L=0.186U  W=1.14U   
+  PD=1.069U
M7      U9_drain A1      U8_source VDD     P   L=0.18U  W=1.51U   
+  PS=1.030U PD=1.030U
M8      U8_source U10_gate VDD     VDD     P   L=0.18U  W=1.51U   
+  PD=1.030U
M9      U4_drain A2      VDD     VDD     P   L=0.18U  W=1.51U   
+  PD=1.030U
M10     U9_drain U9_gate U4_drain VDD     P   L=0.18U  W=1.51U   
+  PS=1.030U PD=1.030U
M11     Z       U195_gate VDD     VDD     P   L=0.182U  W=14.34U   
+  PD=1.603U
M12     U195_gate U9_drain VDD     VDD     P   L=0.183U  W=3.2U   
+  PD=1.603U
M13     U9_gate A1      VSS     VSS     N   L=0.18U  W=0.42U  
M14     U9_gate A1      VDD     VDD     P   L=0.18U  W=1.15U  
M15     U10_gate A2      VSS     VSS     N   L=0.18U  W=0.42U  
M16     U10_gate A2      VDD     VDD     P   L=0.186U  W=1.19U  

.ENDS xr02d7

.SUBCKT xr02da Z  A1 A2 VDD VSS
M1      U9_drain U9_gate U9_source VSS     N   L=0.18U  W=0.54U   
+  PS=.745U PD=.697U
M2      U9_source U10_gate VSS     VSS     N   L=0.18U  W=0.54U   
+  PD=.745U
M3      U63_drain A2      VSS     VSS     N   L=0.18U  W=0.54U   
+  PD=.613U
M4      U9_drain A1      U63_drain VSS     N   L=0.18U  W=0.54U   
+  PS=.613U PD=.697U
M5      Z       U195_gate VSS     VSS     N   L=0.183U  W=7.09U   
+  PD=1.069U
M6      U195_gate U9_drain VSS     VSS     N   L=0.18U  W=1.43U   
+  PD=1.069U
M7      U9_drain A1      U8_source VDD     P   L=0.18U  W=1.51U   
+  PS=1.030U PD=1.030U
M8      U8_source U10_gate VDD     VDD     P   L=0.18U  W=1.51U   
+  PD=1.030U
M9      U4_drain A2      VDD     VDD     P   L=0.18U  W=1.51U   
+  PD=1.030U
M10     U9_drain U9_gate U4_drain VDD     P   L=0.18U  W=1.51U   
+  PS=1.030U PD=1.030U
M11     Z       U195_gate VDD     VDD     P   L=0.182U  W=20.28U   
+  PD=1.603U
M12     U195_gate U9_drain VDD     VDD     P   L=0.183U  W=3.82U   
+  PD=1.603U
M13     U9_gate A1      VSS     VSS     N   L=0.18U  W=0.42U  
M14     U9_gate A1      VDD     VDD     P   L=0.18U  W=1.15U  
M15     U10_gate A2      VSS     VSS     N   L=0.18U  W=0.42U  
M16     U10_gate A2      VDD     VDD     P   L=0.18U  W=1.19U  

.ENDS xr02da

.SUBCKT xr03d7 Z  A1 A2 A3 VDD VSS
M1      u12_out K       VSS     VSS     N   L=0.18U  W=0.55U  
M2      u12_out K       VDD     VDD     P   L=0.18U  W=1.51U  
M3      u19_G   u19_GB  VSS     VSS     N   L=0.18U  W=0.42U  
M4      u19_G   u19_GB  VDD     VDD     P   L=0.187U  W=1.08U  
M5      u10_G   A2      VSS     VSS     N   L=0.18U  W=0.42U  
M6      u10_G   A2      VDD     VDD     P   L=0.187U  W=1.15U  
M7      D       A3      VSS     VSS     N   L=0.18U  W=0.6U  
M8      D       A3      VDD     VDD     P   L=0.18U  W=1.59U  
M9      u11_S   D       VSS     VSS     N   L=0.18U  W=0.6U  
M10     u11_S   D       VDD     VDD     P   L=0.18U  W=1.51U  
M11     K       A1      VSS     VSS     N   L=0.18U  W=0.55U  
M12     K       A1      VDD     VDD     P   L=0.185U  W=1.55U  
M13     K       u19_GB  u19_D   VDD     P   L=0.18U  W=1.55U  
M14     K       u19_G   u19_D   VSS     N   L=0.18U  W=0.55U  
M15     D       A2      u19_GB  VDD     P   L=0.18U  W=1.59U  
M16     D       u10_G   u19_GB  VSS     N   L=0.18U  W=0.6U  
M17     u11_S   u10_G   u19_GB  VDD     P   L=0.185U  W=1.51U  
M18     u11_S   A2      u19_GB  VSS     N   L=0.18U  W=0.66U  
M19     u12_out u19_G   u19_D   VDD     P   L=0.185U  W=1.51U  
M20     u12_out u19_GB  u19_D   VSS     N   L=0.18U  W=0.55U  
M21     Z       U198_gate VSS     VSS     N   L=0.18U  W=5.07U   
+  PD=1.284U
M22     U198_gate u19_D   VSS     VSS     N   L=0.187U  W=1.15U   
+  PD=1.284U
M23     Z       U198_gate VDD     VDD     P   L=0.182U  W=14.34U   
+  PD=1.484U
M24     U198_gate u19_D   VDD     VDD     P   L=0.1825U  W=3.25U   
+  PD=1.484U

.ENDS xr03d7

.SUBCKT xr03da Z  A1 A2 A3 VDD VSS
M1      u12_out K       VSS     VSS     N   L=0.18U  W=0.58U  
M2      u12_out K       VDD     VDD     P   L=0.185U  W=1.51U  
M3      u19_G   u19_GB  VSS     VSS     N   L=0.18U  W=0.42U  
M4      u19_G   u19_GB  VDD     VDD     P   L=0.18U  W=1.15U  
M5      u10_G   A2      VSS     VSS     N   L=0.18U  W=0.42U  
M6      u10_G   A2      VDD     VDD     P   L=0.186U  W=1.19U  
M7      D       A3      VSS     VSS     N   L=0.18U  W=0.59U  
M8      D       A3      VDD     VDD     P   L=0.18U  W=1.59U  
M9      u11_S   D       VSS     VSS     N   L=0.18U  W=0.59U  
M10     u11_S   D       VDD     VDD     P   L=0.185U  W=1.51U  
M11     K       A1      VSS     VSS     N   L=0.18U  W=0.55U  
M12     K       A1      VDD     VDD     P   L=0.185U  W=1.55U  
M13     K       u19_GB  u19_D   VDD     P   L=0.18U  W=1.55U  
M14     K       u19_G   u19_D   VSS     N   L=0.18U  W=0.55U  
M15     D       A2      u19_GB  VDD     P   L=0.18U  W=1.55U  
M16     D       u10_G   u19_GB  VSS     N   L=0.18U  W=0.59U  
M17     u11_S   u10_G   u19_GB  VDD     P   L=0.18U  W=1.51U  
M18     u11_S   A2      u19_GB  VSS     N   L=0.18U  W=0.66U  
M19     u12_out u19_G   u19_D   VDD     P   L=0.18U  W=1.51U  
M20     u12_out u19_GB  u19_D   VSS     N   L=0.18U  W=0.55U  
M21     Z       U198_gate VSS     VSS     N   L=0.183U  W=7.09U   
+  PD=1.284U
M22     U198_gate u19_D   VSS     VSS     N   L=0.18U  W=1.43U   
+  PD=1.284U
M23     Z       U198_gate VDD     VDD     P   L=0.18225U  W=20.37U   
+  PD=1.484U
M24     U198_gate u19_D   VDD     VDD     P   L=0.183U  W=3.88U   
+  PD=1.484U

.ENDS xr03da

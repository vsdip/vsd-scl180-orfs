

VERSION 5.4 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 1000  ;
    TIME NANOSECONDS 1  ;
    CAPACITANCE PICOFARADS 1  ;
    RESISTANCE OHMS 1  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;
SITE CoreSite
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE 0.560 BY 5.600 ;
END CoreSite

MACRO xr03da
    CLASS CORE ;
    FOREIGN xr03da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.386  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.200 1.990 4.440 3.160 ;
        RECT  3.980 1.990 4.440 2.480 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.298  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.660 1.250 3.110 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.392  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.840 2.010 1.620 2.410 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.677  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.470 1.180 14.990 2.980 ;
        RECT  11.380 1.210 14.990 2.980 ;
        RECT  12.440 1.210 12.940 4.330 ;
        RECT  10.010 2.570 12.940 3.070 ;
        RECT  10.120 1.210 14.990 1.710 ;
        RECT  10.120 1.200 10.520 1.710 ;
        RECT  10.010 2.570 10.510 4.330 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.120 5.600 ;
        RECT  14.560 4.620 14.980 5.600 ;
        RECT  13.270 3.210 13.510 5.600 ;
        RECT  12.060 4.590 12.460 5.600 ;
        RECT  10.750 3.300 11.150 5.600 ;
        RECT  9.630 4.590 10.030 5.600 ;
        RECT  8.320 4.620 8.720 5.600 ;
        RECT  6.700 4.610 7.100 5.600 ;
        RECT  3.680 4.620 4.080 5.600 ;
        RECT  0.750 4.620 1.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.120 0.740 ;
        RECT  13.620 0.000 14.020 0.980 ;
        RECT  12.240 0.000 12.640 0.980 ;
        RECT  10.860 0.000 11.260 0.980 ;
        RECT  9.480 0.000 9.880 0.980 ;
        RECT  7.940 0.000 8.350 0.980 ;
        RECT  6.660 0.000 7.100 1.260 ;
        RECT  3.220 0.000 3.620 0.980 ;
        RECT  0.500 0.000 0.900 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.140 0.980 2.270 1.220 ;
        RECT  1.140 0.980 1.380 1.760 ;
        RECT  0.140 1.480 1.380 1.760 ;
        RECT  0.140 1.480 0.550 1.880 ;
        RECT  0.140 1.480 0.470 2.060 ;
        RECT  0.140 1.480 0.380 3.610 ;
        RECT  0.230 3.360 0.470 4.060 ;
        RECT  3.010 1.720 3.600 1.960 ;
        RECT  3.010 1.720 3.250 3.900 ;
        RECT  3.010 3.480 3.470 3.900 ;
        RECT  1.620 1.510 2.170 1.750 ;
        RECT  1.930 1.510 2.170 2.940 ;
        RECT  1.650 2.700 2.170 2.940 ;
        RECT  3.500 2.200 3.740 3.230 ;
        RECT  1.650 2.700 1.890 4.380 ;
        RECT  3.720 2.990 3.960 4.380 ;
        RECT  1.650 4.140 3.960 4.380 ;
        RECT  4.060 0.990 6.010 1.230 ;
        RECT  4.060 0.990 4.300 1.480 ;
        RECT  2.530 1.240 4.300 1.480 ;
        RECT  2.530 1.240 2.770 2.490 ;
        RECT  2.410 2.250 2.650 3.650 ;
        RECT  6.040 1.980 6.570 2.390 ;
        RECT  6.040 1.980 6.280 3.750 ;
        RECT  4.680 1.470 6.470 1.710 ;
        RECT  6.230 1.500 7.110 1.740 ;
        RECT  4.680 1.470 4.930 2.530 ;
        RECT  6.860 1.500 7.110 3.230 ;
        RECT  6.540 2.820 7.110 3.230 ;
        RECT  4.760 2.270 5.000 4.040 ;
        RECT  4.420 3.640 5.000 4.040 ;
        RECT  7.550 1.220 8.070 1.640 ;
        RECT  7.550 1.220 7.790 3.820 ;
        RECT  5.300 1.950 5.800 2.360 ;
        RECT  8.030 2.530 8.440 2.930 ;
        RECT  5.300 1.950 5.540 4.350 ;
        RECT  8.110 2.530 8.350 4.350 ;
        RECT  5.300 4.110 8.350 4.350 ;
        RECT  8.740 1.280 9.440 1.680 ;
        RECT  9.070 1.940 11.150 2.340 ;
        RECT  9.070 1.280 9.440 4.200 ;
        RECT  8.890 3.790 9.440 4.200 ;
    END
END xr03da

MACRO xr03d7
    CLASS CORE ;
    FOREIGN xr03d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.386  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.580 4.420 3.200 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.290  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.310 1.900 0.710 2.300 ;
        RECT  0.120 2.020 0.500 2.460 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.394  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.670 1.060 3.580 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.960  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.880 2.660 13.320 2.900 ;
        RECT  12.900 1.230 13.320 2.900 ;
        RECT  9.340 1.230 13.320 1.470 ;
        RECT  10.880 2.660 11.120 4.340 ;
        RECT  9.490 3.520 11.120 3.760 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 13.440 5.600 ;
        RECT  12.700 4.100 13.100 5.600 ;
        RECT  11.360 3.260 11.760 5.600 ;
        RECT  10.240 4.620 10.640 5.600 ;
        RECT  8.940 4.620 9.340 5.600 ;
        RECT  7.580 4.620 7.980 5.600 ;
        RECT  6.280 4.400 6.680 5.600 ;
        RECT  3.600 4.590 4.000 5.600 ;
        RECT  0.740 4.400 1.140 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 13.440 0.740 ;
        RECT  11.580 0.000 11.980 0.990 ;
        RECT  10.080 0.000 10.480 0.990 ;
        RECT  8.600 0.000 9.000 0.980 ;
        RECT  6.690 0.000 6.930 2.270 ;
        RECT  3.130 0.000 3.530 0.890 ;
        RECT  0.420 0.000 0.820 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.060 0.980 2.260 1.220 ;
        RECT  0.950 1.130 1.290 1.370 ;
        RECT  0.150 1.410 1.190 1.650 ;
        RECT  0.950 1.130 1.190 2.430 ;
        RECT  0.950 2.190 1.540 2.430 ;
        RECT  1.300 2.190 1.540 4.060 ;
        RECT  0.150 3.820 1.540 4.060 ;
        RECT  3.080 1.630 3.320 2.170 ;
        RECT  2.910 1.940 3.150 3.510 ;
        RECT  1.510 1.470 2.010 1.950 ;
        RECT  1.710 1.950 2.020 2.020 ;
        RECT  1.780 1.950 2.020 2.380 ;
        RECT  3.390 2.400 3.630 3.980 ;
        RECT  2.970 3.750 3.570 3.990 ;
        RECT  1.800 2.210 2.040 4.620 ;
        RECT  2.970 3.750 3.210 4.620 ;
        RECT  1.470 4.380 3.210 4.620 ;
        RECT  3.780 0.980 5.750 1.220 ;
        RECT  2.500 1.130 4.020 1.370 ;
        RECT  2.500 1.130 2.740 1.770 ;
        RECT  2.250 1.460 2.650 1.860 ;
        RECT  2.310 1.460 2.650 1.920 ;
        RECT  2.310 1.460 2.550 4.140 ;
        RECT  5.950 1.940 6.190 3.340 ;
        RECT  5.620 3.070 6.190 3.340 ;
        RECT  5.620 3.070 5.860 3.690 ;
        RECT  6.140 1.130 6.380 1.700 ;
        RECT  4.370 1.460 6.380 1.700 ;
        RECT  4.370 1.460 4.770 2.320 ;
        RECT  4.660 2.070 4.900 3.850 ;
        RECT  4.170 3.610 4.900 3.850 ;
        RECT  7.430 0.980 7.860 1.380 ;
        RECT  7.430 0.980 7.670 2.750 ;
        RECT  6.710 2.510 7.670 2.750 ;
        RECT  6.710 2.510 6.950 3.680 ;
        RECT  6.710 3.440 7.280 3.680 ;
        RECT  5.210 1.940 5.450 2.720 ;
        RECT  7.900 2.920 8.300 3.320 ;
        RECT  7.580 3.000 8.300 3.320 ;
        RECT  5.940 3.920 7.820 4.160 ;
        RECT  7.580 3.000 7.820 4.160 ;
        RECT  5.140 3.930 6.010 4.170 ;
        RECT  5.140 2.400 5.380 4.610 ;
        RECT  4.910 4.210 5.380 4.610 ;
        RECT  8.100 1.240 8.340 2.260 ;
        RECT  8.100 1.860 12.640 2.260 ;
        RECT  8.630 1.860 8.910 3.850 ;
        RECT  8.220 3.610 8.910 3.850 ;
        RECT  8.220 3.610 8.480 4.370 ;
    END
END xr03d7

MACRO xr03d4
    CLASS CORE ;
    FOREIGN xr03d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.330 2.830 6.100 3.070 ;
        RECT  5.640 2.580 6.100 3.070 ;
        RECT  5.640 1.630 5.880 3.070 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.311  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.030 3.020 ;
        RECT  0.620 2.020 1.000 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.329  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.270 2.020 1.620 2.630 ;
        RECT  1.240 2.020 1.620 2.460 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.070 3.360 10.900 3.600 ;
        RECT  8.880 1.630 10.670 1.870 ;
        RECT  9.580 1.630 10.020 3.600 ;
        RECT  8.880 1.630 10.020 1.930 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  9.690 4.620 10.090 5.600 ;
        RECT  8.140 4.610 8.540 5.600 ;
        RECT  5.550 4.400 5.790 5.600 ;
        RECT  4.230 4.270 4.470 5.600 ;
        RECT  1.150 3.770 1.390 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  9.610 0.000 9.850 1.190 ;
        RECT  8.110 0.000 8.510 0.890 ;
        RECT  5.380 0.000 5.620 1.200 ;
        RECT  3.880 0.000 4.280 0.890 ;
        RECT  0.970 0.000 1.210 1.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.460 0.550 1.780 ;
        RECT  0.120 1.460 0.360 3.590 ;
        RECT  0.120 3.270 0.730 3.590 ;
        RECT  0.490 3.270 0.730 4.620 ;
        RECT  0.140 4.380 0.730 4.620 ;
        RECT  3.190 1.490 3.550 3.650 ;
        RECT  1.630 1.460 2.100 1.780 ;
        RECT  1.860 1.460 2.100 4.620 ;
        RECT  1.830 2.870 2.100 4.620 ;
        RECT  1.830 4.380 3.870 4.620 ;
        RECT  2.450 1.490 2.690 2.160 ;
        RECT  3.790 2.600 4.560 2.840 ;
        RECT  2.570 1.950 2.810 4.130 ;
        RECT  3.790 2.600 4.030 4.130 ;
        RECT  2.570 3.890 4.030 4.130 ;
        RECT  4.470 1.570 5.090 1.810 ;
        RECT  4.850 2.070 5.240 2.470 ;
        RECT  4.850 1.570 5.090 3.650 ;
        RECT  7.440 1.610 7.920 1.930 ;
        RECT  7.440 1.610 7.680 3.680 ;
        RECT  7.440 3.360 7.920 3.680 ;
        RECT  6.040 1.130 8.400 1.370 ;
        RECT  6.040 1.100 6.580 1.420 ;
        RECT  8.160 1.130 8.400 2.540 ;
        RECT  7.920 2.220 8.400 2.540 ;
        RECT  6.340 1.100 6.580 3.680 ;
        RECT  6.040 3.360 6.580 3.680 ;
        RECT  8.340 2.830 8.920 3.070 ;
        RECT  6.860 1.610 7.100 4.160 ;
        RECT  8.340 2.830 8.580 4.160 ;
        RECT  6.860 3.920 8.580 4.160 ;
    END
END xr03d4

MACRO xr03d2
    CLASS CORE ;
    FOREIGN xr03d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.330 2.830 6.100 3.070 ;
        RECT  5.640 2.580 6.100 3.070 ;
        RECT  5.640 1.630 5.880 3.070 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.311  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.030 3.020 ;
        RECT  0.620 2.020 1.000 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.329  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.270 2.020 1.620 2.630 ;
        RECT  1.240 2.020 1.620 2.460 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.202  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.940 3.360 9.460 3.680 ;
        RECT  9.160 2.020 9.460 3.680 ;
        RECT  8.960 1.610 9.200 2.460 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  9.610 4.300 9.850 5.600 ;
        RECT  8.220 4.400 8.460 5.600 ;
        RECT  5.550 4.400 5.790 5.600 ;
        RECT  4.240 4.250 4.480 5.600 ;
        RECT  1.150 3.770 1.390 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  9.610 0.000 9.850 1.380 ;
        RECT  8.110 0.000 8.510 0.890 ;
        RECT  5.380 0.000 5.620 1.200 ;
        RECT  3.880 0.000 4.280 1.030 ;
        RECT  0.970 0.000 1.210 1.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.460 0.550 1.780 ;
        RECT  0.120 1.460 0.360 3.590 ;
        RECT  0.120 3.270 0.730 3.590 ;
        RECT  0.490 3.270 0.730 4.620 ;
        RECT  0.140 4.380 0.730 4.620 ;
        RECT  3.190 1.490 3.550 3.650 ;
        RECT  1.630 1.460 2.100 1.780 ;
        RECT  1.860 1.460 2.100 4.620 ;
        RECT  1.830 2.870 2.100 4.620 ;
        RECT  1.830 4.380 3.870 4.620 ;
        RECT  2.450 1.490 2.690 2.160 ;
        RECT  3.790 2.760 4.560 3.000 ;
        RECT  2.570 1.950 2.810 4.130 ;
        RECT  3.790 2.760 4.030 4.130 ;
        RECT  2.570 3.890 4.030 4.130 ;
        RECT  4.470 1.570 5.090 1.810 ;
        RECT  4.850 2.070 5.240 2.470 ;
        RECT  4.850 1.570 5.090 3.650 ;
        RECT  7.440 1.610 7.920 1.930 ;
        RECT  7.440 1.610 7.680 3.680 ;
        RECT  7.440 3.360 7.920 3.680 ;
        RECT  6.040 1.130 8.400 1.370 ;
        RECT  6.040 1.100 6.580 1.420 ;
        RECT  8.160 1.130 8.400 2.540 ;
        RECT  7.920 2.220 8.400 2.540 ;
        RECT  6.340 1.100 6.580 3.680 ;
        RECT  6.040 3.360 6.580 3.680 ;
        RECT  8.340 2.830 8.920 3.070 ;
        RECT  6.860 1.610 7.100 4.160 ;
        RECT  8.340 2.830 8.580 4.160 ;
        RECT  6.860 3.920 8.580 4.160 ;
    END
END xr03d2

MACRO xr03d1
    CLASS CORE ;
    FOREIGN xr03d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.330 2.830 6.100 3.070 ;
        RECT  5.640 2.580 6.100 3.070 ;
        RECT  5.640 1.630 5.880 3.070 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.311  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.030 3.020 ;
        RECT  0.620 2.020 1.000 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.329  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.270 2.020 1.620 2.630 ;
        RECT  1.240 2.020 1.620 2.460 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.054  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.820 3.360 9.400 3.600 ;
        RECT  9.160 1.180 9.400 3.600 ;
        RECT  9.020 1.180 9.400 1.900 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  8.190 4.400 8.430 5.600 ;
        RECT  5.550 4.400 5.790 5.600 ;
        RECT  4.250 4.230 4.490 5.600 ;
        RECT  1.150 3.770 1.390 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.210 0.000 8.600 0.890 ;
        RECT  5.470 0.000 5.710 1.200 ;
        RECT  3.930 0.000 4.170 1.750 ;
        RECT  0.970 0.000 1.210 1.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.460 0.550 1.780 ;
        RECT  0.120 1.460 0.360 3.590 ;
        RECT  0.120 3.270 0.730 3.590 ;
        RECT  0.490 3.270 0.730 4.620 ;
        RECT  0.140 4.380 0.730 4.620 ;
        RECT  3.190 1.490 3.550 3.650 ;
        RECT  1.630 1.460 2.100 1.780 ;
        RECT  1.860 1.460 2.100 4.620 ;
        RECT  1.830 2.870 2.100 4.620 ;
        RECT  1.830 4.380 3.870 4.620 ;
        RECT  2.450 1.490 2.690 2.160 ;
        RECT  3.790 2.600 4.560 2.840 ;
        RECT  2.570 1.950 2.810 4.130 ;
        RECT  3.790 2.600 4.030 4.130 ;
        RECT  2.570 3.890 4.030 4.130 ;
        RECT  4.590 1.490 5.090 1.810 ;
        RECT  4.850 2.070 5.240 2.470 ;
        RECT  4.850 1.490 5.090 3.650 ;
        RECT  7.440 1.690 8.010 1.930 ;
        RECT  7.440 1.690 7.680 3.680 ;
        RECT  7.440 3.360 7.920 3.680 ;
        RECT  6.130 1.130 8.540 1.370 ;
        RECT  6.130 1.100 6.580 1.420 ;
        RECT  8.300 1.130 8.540 2.460 ;
        RECT  7.920 2.220 8.540 2.460 ;
        RECT  6.340 1.100 6.580 3.680 ;
        RECT  6.040 3.360 6.580 3.680 ;
        RECT  8.340 2.750 8.920 3.070 ;
        RECT  6.860 1.610 7.190 4.160 ;
        RECT  8.340 2.750 8.580 4.160 ;
        RECT  6.860 3.920 8.580 4.160 ;
    END
END xr03d1

MACRO xr02da
    CLASS CORE ;
    FOREIGN xr02da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.283  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.580 2.580 1.060 3.020 ;
        RECT  0.580 1.980 0.980 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.290  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.410 4.420 3.020 ;
        RECT  3.980 2.090 4.380 3.020 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.347  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.160 1.780 11.610 2.460 ;
        RECT  11.200 1.140 11.610 2.460 ;
        RECT  10.540 1.780 10.940 4.310 ;
        RECT  6.640 2.610 10.940 3.890 ;
        RECT  8.160 1.780 10.940 3.890 ;
        RECT  8.160 1.230 10.220 3.890 ;
        RECT  9.240 1.230 9.640 4.040 ;
        RECT  7.940 2.610 8.340 3.990 ;
        RECT  6.990 1.230 10.220 1.730 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.760 5.600 ;
        RECT  11.200 3.050 11.600 5.600 ;
        RECT  9.980 4.620 10.380 5.600 ;
        RECT  8.680 4.550 9.080 5.600 ;
        RECT  7.380 4.550 7.780 5.600 ;
        RECT  6.080 4.120 6.480 5.600 ;
        RECT  4.780 3.540 5.180 5.600 ;
        RECT  3.180 4.000 3.580 5.600 ;
        RECT  0.750 4.710 1.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.760 0.740 ;
        RECT  10.460 0.000 10.860 1.540 ;
        RECT  9.090 0.000 9.490 0.980 ;
        RECT  7.730 0.000 8.130 0.990 ;
        RECT  6.380 0.000 6.780 0.980 ;
        RECT  4.900 0.000 5.300 1.570 ;
        RECT  3.470 0.000 3.870 0.890 ;
        RECT  0.930 0.000 1.330 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.500 1.830 1.740 ;
        RECT  1.680 1.550 2.770 1.790 ;
        RECT  1.810 1.550 2.050 3.500 ;
        RECT  0.150 3.260 2.050 3.500 ;
        RECT  3.490 1.610 4.420 1.850 ;
        RECT  3.490 1.610 3.730 2.920 ;
        RECT  2.930 2.590 3.730 2.920 ;
        RECT  2.930 2.590 3.330 3.760 ;
        RECT  2.930 3.520 4.240 3.760 ;
        RECT  4.000 3.520 4.240 4.390 ;
        RECT  2.020 0.980 3.240 1.220 ;
        RECT  4.210 0.990 4.610 1.370 ;
        RECT  3.010 1.130 4.610 1.370 ;
        RECT  3.010 1.130 3.250 2.320 ;
        RECT  2.290 2.080 3.250 2.320 ;
        RECT  2.290 2.080 2.530 4.000 ;
        RECT  1.980 3.760 2.530 4.000 ;
        RECT  5.640 1.250 6.400 1.650 ;
        RECT  6.000 1.980 7.910 2.380 ;
        RECT  6.000 1.250 6.400 3.130 ;
        RECT  5.340 2.730 6.400 3.130 ;
    END
END xr02da

MACRO xr02d7
    CLASS CORE ;
    FOREIGN xr02d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.283  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.980 0.800 2.380 ;
        RECT  0.120 1.980 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.298  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.340 2.560 4.980 3.020 ;
        RECT  3.960 2.490 4.580 2.730 ;
        RECT  3.960 2.170 4.200 2.730 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.620 1.250 9.850 1.650 ;
        RECT  9.450 0.980 9.850 1.650 ;
        RECT  8.960 2.580 9.460 3.020 ;
        RECT  6.540 2.570 9.420 2.970 ;
        RECT  9.020 1.250 9.420 3.020 ;
        RECT  8.960 2.570 9.360 3.800 ;
        RECT  7.660 2.570 8.060 4.340 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  9.530 4.620 9.930 5.600 ;
        RECT  8.220 4.620 8.620 5.600 ;
        RECT  7.180 3.260 7.420 5.600 ;
        RECT  5.800 3.950 6.200 5.600 ;
        RECT  4.490 3.950 4.890 5.600 ;
        RECT  3.290 3.520 3.530 5.600 ;
        RECT  0.570 4.710 0.970 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  8.680 0.000 9.080 0.980 ;
        RECT  7.360 0.000 7.760 0.980 ;
        RECT  5.880 0.000 6.280 0.990 ;
        RECT  3.500 0.000 3.900 0.890 ;
        RECT  0.930 0.000 1.330 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.500 1.830 1.740 ;
        RECT  1.750 1.510 2.760 1.750 ;
        RECT  1.800 1.510 2.040 3.500 ;
        RECT  0.150 3.260 2.040 3.500 ;
        RECT  3.480 1.610 4.660 1.850 ;
        RECT  3.480 1.610 3.720 2.710 ;
        RECT  2.940 2.470 3.720 2.710 ;
        RECT  3.260 2.470 3.500 3.280 ;
        RECT  3.260 3.040 4.100 3.280 ;
        RECT  3.860 3.040 4.100 4.610 ;
        RECT  2.010 0.980 3.240 1.220 ;
        RECT  3.000 1.130 5.140 1.370 ;
        RECT  4.900 1.130 5.140 2.290 ;
        RECT  3.000 0.980 3.240 2.230 ;
        RECT  2.330 1.990 3.240 2.230 ;
        RECT  4.900 2.050 5.630 2.290 ;
        RECT  5.390 2.050 5.630 2.680 ;
        RECT  2.330 1.990 2.570 4.000 ;
        RECT  2.000 3.760 2.570 4.000 ;
        RECT  5.380 1.250 5.620 1.810 ;
        RECT  5.380 1.570 6.210 1.810 ;
        RECT  5.910 1.570 6.210 2.330 ;
        RECT  5.910 1.930 8.670 2.330 ;
        RECT  5.910 1.570 6.150 3.520 ;
        RECT  5.060 3.280 6.150 3.520 ;
    END
END xr02d7

MACRO xr02d4
    CLASS CORE ;
    FOREIGN xr02d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.263  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.700 2.740 4.520 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.346  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 1.620 2.920 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.068  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.780 1.750 6.550 1.990 ;
        RECT  4.610 3.130 6.330 3.370 ;
        RECT  5.100 1.750 5.540 3.370 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.200 4.620 5.600 5.600 ;
        RECT  3.820 3.610 4.060 5.600 ;
        RECT  1.020 3.990 1.260 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.460 0.000 5.860 0.980 ;
        RECT  4.120 0.000 4.360 1.560 ;
        RECT  1.060 0.000 1.460 1.050 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 1.290 2.630 1.530 ;
        RECT  2.390 1.290 2.630 2.050 ;
        RECT  0.200 1.290 0.610 2.170 ;
        RECT  0.200 1.290 0.440 4.310 ;
        RECT  0.200 3.990 0.600 4.310 ;
        RECT  1.860 2.600 3.840 2.840 ;
        RECT  1.860 1.770 2.100 3.400 ;
        RECT  0.690 3.160 2.100 3.400 ;
        RECT  2.920 1.410 3.160 2.280 ;
        RECT  2.920 2.040 4.320 2.280 ;
        RECT  4.080 2.520 4.630 2.760 ;
        RECT  4.080 2.040 4.320 3.370 ;
        RECT  2.490 3.130 4.320 3.370 ;
    END
END xr02d4

MACRO xr02d2
    CLASS CORE ;
    FOREIGN xr02d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.263  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.700 2.740 4.620 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.346  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 1.620 2.920 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.332  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.580 5.540 3.020 ;
        RECT  4.720 3.750 5.340 3.990 ;
        RECT  5.100 1.750 5.340 3.990 ;
        RECT  4.780 1.750 5.340 1.990 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.650 4.050 5.890 5.600 ;
        RECT  3.950 3.610 4.190 5.600 ;
        RECT  1.020 3.990 1.260 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.590 0.000 5.830 1.560 ;
        RECT  4.120 0.000 4.360 1.560 ;
        RECT  1.060 0.000 1.460 1.050 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 1.290 2.630 1.530 ;
        RECT  2.390 1.290 2.630 2.050 ;
        RECT  0.200 1.290 0.610 2.170 ;
        RECT  0.200 1.290 0.440 4.310 ;
        RECT  0.200 3.990 0.600 4.310 ;
        RECT  1.860 2.600 3.950 2.840 ;
        RECT  1.860 1.770 2.100 3.400 ;
        RECT  0.690 3.160 2.100 3.400 ;
        RECT  2.920 1.410 3.160 2.280 ;
        RECT  2.920 2.040 4.430 2.280 ;
        RECT  4.190 2.200 4.630 2.600 ;
        RECT  4.190 2.040 4.430 3.370 ;
        RECT  2.490 3.130 4.430 3.370 ;
    END
END xr02d2

MACRO xr02d1
    CLASS CORE ;
    FOREIGN xr02d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.263  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.700 2.740 4.620 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.346  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 1.620 2.920 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.046  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.640 3.830 5.480 4.070 ;
        RECT  5.100 1.670 5.480 4.070 ;
        RECT  4.880 1.670 5.480 2.070 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  3.950 3.610 4.190 5.600 ;
        RECT  1.020 3.990 1.260 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.210 0.000 4.450 1.560 ;
        RECT  1.060 0.000 1.460 1.050 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 1.290 2.630 1.530 ;
        RECT  2.390 1.290 2.630 2.050 ;
        RECT  0.200 1.290 0.610 2.170 ;
        RECT  0.200 1.290 0.440 4.310 ;
        RECT  0.200 3.990 0.600 4.310 ;
        RECT  1.860 2.600 4.010 2.840 ;
        RECT  1.860 1.770 2.100 3.400 ;
        RECT  0.690 3.160 2.100 3.400 ;
        RECT  3.010 1.410 3.250 2.280 ;
        RECT  3.010 2.040 4.640 2.280 ;
        RECT  4.400 2.040 4.640 3.370 ;
        RECT  2.490 3.130 4.640 3.370 ;
    END
END xr02d1

MACRO xn02da
    CLASS CORE ;
    FOREIGN xn02da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.150 3.900 3.580 ;
        RECT  3.660 2.600 3.900 3.580 ;
        RECT  3.440 3.140 3.900 3.580 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.648  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.810 2.920 ;
        RECT  0.120 2.580 0.510 3.020 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.569  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.290 1.240 11.640 3.720 ;
        RECT  6.400 2.580 11.640 2.940 ;
        RECT  8.460 1.240 11.640 2.940 ;
        RECT  8.820 1.240 9.060 4.340 ;
        RECT  7.170 1.240 11.640 1.700 ;
        RECT  6.400 2.580 6.640 4.350 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.760 5.600 ;
        RECT  10.640 4.010 11.040 5.600 ;
        RECT  9.380 3.240 9.620 5.600 ;
        RECT  8.180 4.620 8.580 5.600 ;
        RECT  6.960 3.250 7.200 5.600 ;
        RECT  5.740 4.620 6.140 5.600 ;
        RECT  4.430 4.230 4.830 5.600 ;
        RECT  3.020 4.610 3.420 5.600 ;
        RECT  0.630 4.710 1.030 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.760 0.740 ;
        RECT  10.860 0.000 11.260 0.920 ;
        RECT  9.420 0.000 9.820 0.900 ;
        RECT  7.920 0.000 8.320 0.900 ;
        RECT  6.480 0.000 6.880 0.900 ;
        RECT  5.120 0.000 5.360 1.660 ;
        RECT  3.580 0.000 3.820 0.890 ;
        RECT  0.830 0.000 1.070 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.610 1.350 1.860 ;
        RECT  1.110 2.060 1.490 2.470 ;
        RECT  1.080 2.100 1.490 2.470 ;
        RECT  2.880 2.620 3.280 2.940 ;
        RECT  2.880 2.620 3.180 3.410 ;
        RECT  2.580 3.170 3.180 3.410 ;
        RECT  0.150 3.260 1.350 3.500 ;
        RECT  1.110 1.610 1.350 4.060 ;
        RECT  2.580 3.170 2.820 4.060 ;
        RECT  1.110 3.820 2.820 4.060 ;
        RECT  0.160 0.980 0.560 1.370 ;
        RECT  1.300 0.980 3.350 1.220 ;
        RECT  0.160 1.130 1.540 1.370 ;
        RECT  4.070 1.610 4.630 1.850 ;
        RECT  4.390 1.610 4.630 2.350 ;
        RECT  2.280 2.110 4.630 2.350 ;
        RECT  2.280 2.110 2.520 2.930 ;
        RECT  4.070 3.750 4.380 3.990 ;
        RECT  4.140 2.110 4.380 3.990 ;
        RECT  3.690 3.820 4.260 4.060 ;
        RECT  4.070 0.980 4.880 1.220 ;
        RECT  3.590 1.130 4.310 1.370 ;
        RECT  3.590 1.130 3.830 1.760 ;
        RECT  1.730 1.520 3.830 1.760 ;
        RECT  1.730 1.520 1.970 3.500 ;
        RECT  1.730 3.260 2.320 3.500 ;
        RECT  5.750 1.240 6.150 2.340 ;
        RECT  5.080 1.930 6.150 2.340 ;
        RECT  5.080 1.940 8.220 2.340 ;
        RECT  5.080 1.930 5.480 3.900 ;
    END
END xn02da

MACRO xn02d7
    CLASS CORE ;
    FOREIGN xn02d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.140 3.900 3.580 ;
        RECT  3.660 2.600 3.900 3.580 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.648  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.810 2.920 ;
        RECT  0.120 2.520 0.510 3.020 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.519  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.370 2.740 9.960 2.980 ;
        RECT  9.440 1.410 9.960 2.980 ;
        RECT  6.980 1.410 9.960 1.650 ;
        RECT  7.670 2.740 7.910 4.550 ;
        RECT  6.370 2.740 6.610 4.350 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  9.480 4.430 9.880 5.600 ;
        RECT  8.230 3.470 8.470 5.600 ;
        RECT  6.930 3.220 7.170 5.600 ;
        RECT  5.730 4.620 6.130 5.600 ;
        RECT  4.490 4.200 4.730 5.600 ;
        RECT  3.020 4.620 3.420 5.600 ;
        RECT  0.630 4.710 1.030 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  9.530 0.000 9.930 1.010 ;
        RECT  7.740 0.000 8.150 1.010 ;
        RECT  6.410 0.000 6.810 1.010 ;
        RECT  4.870 1.500 5.450 1.740 ;
        RECT  5.210 0.000 5.450 1.740 ;
        RECT  3.580 0.000 3.820 0.890 ;
        RECT  0.830 0.000 1.070 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.610 1.350 1.860 ;
        RECT  1.110 2.060 1.490 2.470 ;
        RECT  1.080 2.100 1.490 2.470 ;
        RECT  2.880 2.620 3.280 2.940 ;
        RECT  2.880 2.620 3.180 3.410 ;
        RECT  2.580 3.170 3.180 3.410 ;
        RECT  0.150 3.260 1.350 3.500 ;
        RECT  1.110 1.610 1.350 4.060 ;
        RECT  2.580 3.170 2.820 4.060 ;
        RECT  1.110 3.820 2.820 4.060 ;
        RECT  0.160 0.980 0.560 1.370 ;
        RECT  1.310 0.980 3.350 1.220 ;
        RECT  0.160 1.130 1.550 1.370 ;
        RECT  4.070 1.610 4.630 1.850 ;
        RECT  4.390 1.610 4.630 2.350 ;
        RECT  2.280 2.110 4.630 2.350 ;
        RECT  2.280 2.110 2.520 2.930 ;
        RECT  4.080 3.760 4.380 3.970 ;
        RECT  4.140 2.110 4.380 3.970 ;
        RECT  3.690 3.820 4.270 4.060 ;
        RECT  4.070 0.980 4.880 1.220 ;
        RECT  3.590 1.130 4.310 1.370 ;
        RECT  3.590 1.130 3.830 1.760 ;
        RECT  1.780 1.520 3.830 1.760 ;
        RECT  1.780 1.520 2.020 2.410 ;
        RECT  1.730 2.170 1.970 3.500 ;
        RECT  1.730 3.260 2.320 3.500 ;
        RECT  5.720 1.290 5.960 2.400 ;
        RECT  5.050 2.160 8.720 2.400 ;
        RECT  5.050 2.160 5.290 3.980 ;
    END
END xn02d7

MACRO xn02d4
    CLASS CORE ;
    FOREIGN xn02d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.532  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.240 0.810 2.480 ;
        RECT  0.120 2.240 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.020 4.420 2.980 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.695  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.410 3.130 7.120 3.370 ;
        RECT  5.420 1.810 7.120 2.050 ;
        RECT  6.220 1.810 6.660 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.230 4.450 6.470 5.600 ;
        RECT  4.910 4.450 5.150 5.600 ;
        RECT  3.610 4.260 3.850 5.600 ;
        RECT  1.050 4.260 1.290 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.240 0.000 6.480 1.320 ;
        RECT  4.920 0.000 5.160 1.320 ;
        RECT  3.450 0.000 3.690 1.300 ;
        RECT  0.940 0.000 1.340 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.300 1.780 ;
        RECT  1.060 2.340 2.660 2.580 ;
        RECT  1.060 1.540 1.300 3.560 ;
        RECT  0.310 3.320 1.300 3.560 ;
        RECT  0.310 3.320 0.550 4.450 ;
        RECT  4.220 1.080 4.460 1.780 ;
        RECT  3.380 1.540 4.460 1.780 ;
        RECT  3.380 1.540 3.620 3.500 ;
        RECT  3.380 3.260 4.530 3.500 ;
        RECT  2.140 1.710 3.140 1.950 ;
        RECT  2.900 3.740 5.170 3.980 ;
        RECT  4.930 2.510 5.170 3.980 ;
        RECT  2.900 1.710 3.140 4.100 ;
        RECT  2.330 3.860 3.140 4.100 ;
    END
END xn02d4

MACRO xn02d2
    CLASS CORE ;
    FOREIGN xn02d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.529  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.240 0.810 2.480 ;
        RECT  0.120 2.240 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.020 4.420 2.980 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.162  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.610 3.130 6.100 3.580 ;
        RECT  5.610 1.770 5.850 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  6.230 4.170 6.470 5.600 ;
        RECT  4.880 4.220 5.120 5.600 ;
        RECT  3.790 4.260 4.030 5.600 ;
        RECT  1.230 4.260 1.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  6.170 0.000 6.570 0.940 ;
        RECT  4.870 0.000 5.110 2.170 ;
        RECT  3.480 0.000 3.720 1.300 ;
        RECT  0.920 0.000 1.320 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.300 1.780 ;
        RECT  1.060 2.340 2.660 2.580 ;
        RECT  1.060 1.540 1.300 3.560 ;
        RECT  0.490 3.320 1.300 3.560 ;
        RECT  0.490 3.320 0.730 4.450 ;
        RECT  4.250 1.080 4.490 1.780 ;
        RECT  3.380 1.540 4.490 1.780 ;
        RECT  3.380 1.540 3.620 3.500 ;
        RECT  3.380 3.260 4.710 3.500 ;
        RECT  2.170 1.710 3.140 1.950 ;
        RECT  2.510 3.240 3.140 3.480 ;
        RECT  2.900 1.710 3.140 3.980 ;
        RECT  5.000 2.600 5.240 3.980 ;
        RECT  2.900 3.740 5.240 3.980 ;
    END
END xn02d2

MACRO xn02d1
    CLASS CORE ;
    FOREIGN xn02d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.529  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.240 0.810 2.480 ;
        RECT  0.120 2.240 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.020 4.420 2.980 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.064  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 1.460 6.040 3.450 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.090 4.220 5.330 5.600 ;
        RECT  3.790 4.260 4.030 5.600 ;
        RECT  1.230 4.260 1.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.950 0.000 5.190 1.490 ;
        RECT  3.480 0.000 3.720 1.300 ;
        RECT  0.920 0.000 1.320 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.300 1.780 ;
        RECT  1.060 2.340 2.660 2.580 ;
        RECT  1.060 1.540 1.300 3.560 ;
        RECT  0.490 3.320 1.300 3.560 ;
        RECT  0.490 3.320 0.730 4.450 ;
        RECT  4.250 1.080 4.490 1.780 ;
        RECT  3.380 1.540 4.490 1.780 ;
        RECT  3.380 1.540 3.620 3.500 ;
        RECT  3.380 3.260 4.710 3.500 ;
        RECT  2.170 1.710 3.140 1.950 ;
        RECT  2.510 3.240 3.140 3.480 ;
        RECT  2.900 1.710 3.140 3.980 ;
        RECT  5.180 2.520 5.420 3.980 ;
        RECT  2.900 3.740 5.420 3.980 ;
    END
END xn02d1

MACRO su01d4
    CLASS CORE ;
    FOREIGN su01d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.153  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.150 2.290 7.570 2.530 ;
        RECT  3.540 2.750 5.550 2.990 ;
        RECT  5.150 1.960 5.550 2.990 ;
        RECT  5.100 2.580 5.540 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.328  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.180 2.600 1.420 3.580 ;
        RECT  0.600 2.600 1.420 2.840 ;
        RECT  0.600 2.600 0.840 3.160 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.762  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.740 2.250 4.870 2.490 ;
        RECT  2.300 2.220 3.200 2.460 ;
        RECT  2.300 2.000 2.780 2.460 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.813  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.620 1.340 14.410 1.580 ;
        RECT  14.010 1.180 14.410 1.580 ;
        RECT  12.220 2.690 14.250 2.930 ;
        RECT  14.010 1.180 14.250 2.930 ;
        RECT  13.500 2.580 14.250 2.930 ;
        RECT  13.500 2.580 13.940 3.020 ;
        RECT  13.520 2.580 13.760 4.620 ;
        RECT  12.620 1.180 13.020 1.580 ;
        RECT  12.220 2.690 12.460 4.620 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.035  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.750 1.340 11.540 1.580 ;
        RECT  11.140 1.180 11.540 1.580 ;
        RECT  10.700 2.580 11.360 3.020 ;
        RECT  10.820 2.500 11.360 3.020 ;
        RECT  11.120 1.340 11.360 3.020 ;
        RECT  9.530 2.580 11.360 2.820 ;
        RECT  9.750 1.180 10.150 1.580 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 14.560 5.600 ;
        RECT  14.000 3.530 14.400 5.600 ;
        RECT  12.700 3.520 13.100 5.600 ;
        RECT  11.400 4.620 11.800 5.600 ;
        RECT  10.100 4.620 10.500 5.600 ;
        RECT  7.350 4.650 7.750 5.600 ;
        RECT  6.190 4.650 6.590 5.600 ;
        RECT  3.070 4.340 3.630 4.580 ;
        RECT  3.070 4.340 3.310 5.600 ;
        RECT  0.720 4.120 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 14.560 0.740 ;
        RECT  13.360 0.000 13.760 0.990 ;
        RECT  11.880 0.000 12.280 1.200 ;
        RECT  10.400 0.000 10.800 0.990 ;
        RECT  7.510 0.000 7.910 0.890 ;
        RECT  6.330 0.000 6.730 0.890 ;
        RECT  3.520 0.000 3.920 0.890 ;
        RECT  0.600 0.000 1.000 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.270 0.550 1.670 ;
        RECT  0.120 1.350 1.400 1.670 ;
        RECT  1.160 1.350 1.400 2.350 ;
        RECT  0.120 1.270 0.360 3.820 ;
        RECT  0.120 3.500 0.550 3.820 ;
        RECT  2.480 3.350 4.200 3.590 ;
        RECT  2.750 1.440 4.150 1.680 ;
        RECT  3.910 1.440 4.150 1.960 ;
        RECT  3.910 1.720 4.510 1.960 ;
        RECT  7.520 3.250 8.500 3.490 ;
        RECT  6.760 3.270 8.090 3.510 ;
        RECT  8.280 1.050 8.680 1.550 ;
        RECT  6.920 1.310 8.680 1.550 ;
        RECT  4.640 1.020 6.040 1.260 ;
        RECT  5.800 1.020 6.040 2.030 ;
        RECT  9.100 1.180 9.340 2.330 ;
        RECT  5.800 1.790 9.340 2.030 ;
        RECT  8.910 1.930 10.240 2.330 ;
        RECT  6.230 2.770 9.150 3.010 ;
        RECT  6.230 2.770 6.470 3.700 ;
        RECT  4.500 3.460 6.470 3.700 ;
        RECT  8.910 1.790 9.150 4.110 ;
        RECT  1.660 1.260 2.410 1.500 ;
        RECT  13.030 1.930 13.430 2.330 ;
        RECT  11.650 2.090 13.430 2.330 ;
        RECT  1.660 1.260 1.900 2.900 ;
        RECT  11.650 2.090 11.890 3.800 ;
        RECT  9.390 3.560 11.890 3.800 ;
        RECT  1.900 2.660 2.140 4.530 ;
        RECT  1.900 3.830 4.260 4.070 ;
        RECT  6.950 3.830 8.440 4.070 ;
        RECT  4.020 3.960 7.190 4.200 ;
        RECT  8.200 3.830 8.440 4.620 ;
        RECT  1.900 3.830 2.330 4.530 ;
        RECT  9.390 3.560 9.630 4.620 ;
        RECT  8.200 4.380 9.630 4.620 ;
    END
END su01d4

MACRO su01d2
    CLASS CORE ;
    FOREIGN su01d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.948  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.350 2.680 2.590 ;
        RECT  0.400 2.350 1.060 3.030 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.394  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.160 2.580 8.900 3.190 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.675  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.210 2.020 6.660 3.030 ;
        RECT  4.850 2.120 6.660 2.360 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.231  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.000 3.160 11.700 3.580 ;
        RECT  11.460 1.720 11.700 3.580 ;
        RECT  11.000 1.720 11.700 2.120 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.231  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.580 3.150 10.140 3.580 ;
        RECT  9.900 1.720 10.140 3.580 ;
        RECT  9.700 1.720 10.140 2.120 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.320 5.600 ;
        RECT  11.640 4.290 11.880 5.600 ;
        RECT  10.340 4.310 10.580 5.600 ;
        RECT  8.930 4.710 9.330 5.600 ;
        RECT  7.650 4.710 8.050 5.600 ;
        RECT  4.600 4.710 5.000 5.600 ;
        RECT  2.960 4.040 3.630 4.280 ;
        RECT  2.960 4.040 3.200 5.600 ;
        RECT  0.800 3.960 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.320 0.740 ;
        RECT  11.560 0.000 11.970 1.420 ;
        RECT  10.260 0.000 10.660 1.420 ;
        RECT  7.820 0.000 8.220 0.890 ;
        RECT  4.650 0.000 4.890 1.260 ;
        RECT  3.310 0.000 3.550 1.260 ;
        RECT  0.800 0.000 1.040 1.260 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.300 1.780 3.540 ;
        RECT  1.540 3.300 1.780 4.330 ;
        RECT  1.280 0.980 1.860 1.220 ;
        RECT  1.280 0.980 1.520 1.880 ;
        RECT  0.150 1.640 1.520 1.880 ;
        RECT  3.790 3.080 4.590 3.320 ;
        RECT  4.350 3.080 4.590 3.970 ;
        RECT  4.350 3.730 5.570 3.970 ;
        RECT  3.830 1.580 5.740 1.820 ;
        RECT  7.620 1.750 8.740 1.990 ;
        RECT  7.620 1.750 7.860 3.720 ;
        RECT  7.620 3.480 8.650 3.720 ;
        RECT  6.940 1.130 9.460 1.370 ;
        RECT  6.130 1.420 7.180 1.660 ;
        RECT  9.220 1.130 9.460 2.910 ;
        RECT  9.220 2.510 9.660 2.910 ;
        RECT  6.940 1.130 7.180 3.570 ;
        RECT  5.930 3.330 7.180 3.570 ;
        RECT  2.030 1.740 3.240 1.980 ;
        RECT  3.000 2.600 5.880 2.840 ;
        RECT  10.380 2.600 11.150 2.840 ;
        RECT  5.480 2.600 5.880 3.030 ;
        RECT  2.030 3.240 3.240 3.480 ;
        RECT  3.000 1.740 3.240 3.800 ;
        RECT  3.000 3.560 4.110 3.800 ;
        RECT  10.380 2.600 10.620 4.070 ;
        RECT  9.140 3.830 10.620 4.070 ;
        RECT  3.870 3.560 4.110 4.470 ;
        RECT  9.140 3.830 9.380 4.470 ;
        RECT  3.870 4.230 9.380 4.470 ;
    END
END su01d2

MACRO su01d1
    CLASS CORE ;
    FOREIGN su01d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.948  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.350 2.680 2.590 ;
        RECT  0.400 2.350 1.060 3.030 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.160 3.010 8.820 3.250 ;
        RECT  8.540 2.580 8.820 3.250 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.675  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.210 2.020 6.660 3.030 ;
        RECT  4.850 2.120 6.660 2.360 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.170  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.290 3.320 11.060 3.720 ;
        RECT  10.780 1.770 11.060 3.720 ;
        RECT  10.540 1.770 11.060 2.170 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.113  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.100 1.770 9.570 2.170 ;
        RECT  9.060 3.160 9.380 3.560 ;
        RECT  9.100 1.770 9.380 3.560 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  9.630 4.290 9.870 5.600 ;
        RECT  7.650 4.710 8.050 5.600 ;
        RECT  4.600 4.710 5.000 5.600 ;
        RECT  2.960 4.040 3.630 4.280 ;
        RECT  2.960 4.040 3.200 5.600 ;
        RECT  0.800 3.960 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  9.930 0.000 10.330 1.520 ;
        RECT  7.820 0.000 8.220 0.890 ;
        RECT  4.650 0.000 4.890 1.260 ;
        RECT  3.310 0.000 3.550 1.260 ;
        RECT  0.800 0.000 1.040 1.260 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.300 1.780 3.540 ;
        RECT  1.540 3.300 1.780 4.330 ;
        RECT  1.280 0.980 1.860 1.220 ;
        RECT  1.280 0.980 1.520 1.880 ;
        RECT  0.150 1.640 1.520 1.880 ;
        RECT  3.790 3.080 4.590 3.320 ;
        RECT  4.350 3.080 4.590 3.970 ;
        RECT  4.350 3.730 5.570 3.970 ;
        RECT  3.830 1.580 5.740 1.820 ;
        RECT  8.550 1.670 8.790 2.320 ;
        RECT  7.420 2.080 8.790 2.320 ;
        RECT  7.420 2.080 7.940 2.600 ;
        RECT  7.420 2.080 7.660 3.900 ;
        RECT  7.420 3.660 8.650 3.900 ;
        RECT  8.480 0.980 9.230 1.220 ;
        RECT  6.940 1.130 8.720 1.370 ;
        RECT  6.130 1.420 7.180 1.660 ;
        RECT  6.940 1.130 7.180 3.570 ;
        RECT  5.930 3.330 7.180 3.570 ;
        RECT  2.030 1.740 3.240 1.980 ;
        RECT  3.000 2.600 5.880 2.840 ;
        RECT  9.810 2.710 10.520 2.950 ;
        RECT  5.480 2.600 5.880 3.030 ;
        RECT  2.030 3.240 3.240 3.480 ;
        RECT  3.000 1.740 3.240 3.800 ;
        RECT  3.000 3.560 4.110 3.800 ;
        RECT  9.810 2.710 10.050 4.040 ;
        RECT  9.140 3.800 10.050 4.040 ;
        RECT  3.870 3.560 4.110 4.470 ;
        RECT  9.140 3.800 9.380 4.470 ;
        RECT  3.870 4.230 9.380 4.470 ;
    END
END su01d1

MACRO su01d0
    CLASS CORE ;
    FOREIGN su01d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.948  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.350 2.680 2.590 ;
        RECT  0.400 2.350 1.060 3.030 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.160 3.010 8.820 3.250 ;
        RECT  8.540 2.580 8.820 3.250 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.675  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.210 2.020 6.660 3.030 ;
        RECT  4.850 2.120 6.660 2.360 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.632  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.290 4.020 11.060 4.420 ;
        RECT  10.780 1.770 11.060 4.420 ;
        RECT  10.550 1.770 11.060 2.170 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.863  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.060 1.770 9.570 2.170 ;
        RECT  9.060 1.770 9.380 3.450 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  9.630 4.310 9.870 5.600 ;
        RECT  7.650 4.710 8.050 5.600 ;
        RECT  4.600 4.710 5.000 5.600 ;
        RECT  2.960 4.040 3.630 4.280 ;
        RECT  2.960 4.040 3.200 5.600 ;
        RECT  0.800 3.960 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  9.960 0.000 10.360 0.890 ;
        RECT  7.820 0.000 8.220 0.890 ;
        RECT  4.650 0.000 4.890 1.260 ;
        RECT  3.310 0.000 3.550 1.260 ;
        RECT  0.800 0.000 1.040 1.260 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.300 1.780 3.540 ;
        RECT  1.540 3.300 1.780 4.330 ;
        RECT  1.280 0.980 1.860 1.220 ;
        RECT  1.280 0.980 1.520 1.880 ;
        RECT  0.150 1.640 1.520 1.880 ;
        RECT  3.790 3.080 4.590 3.320 ;
        RECT  4.350 3.080 4.590 3.970 ;
        RECT  4.350 3.730 5.570 3.970 ;
        RECT  3.830 1.580 5.740 1.820 ;
        RECT  8.550 1.670 8.790 2.320 ;
        RECT  7.420 2.080 8.790 2.320 ;
        RECT  7.420 2.080 7.940 2.600 ;
        RECT  7.420 2.080 7.660 3.900 ;
        RECT  7.420 3.660 8.650 3.900 ;
        RECT  6.940 1.130 10.050 1.370 ;
        RECT  6.130 1.420 7.180 1.660 ;
        RECT  9.810 1.130 10.050 2.730 ;
        RECT  9.620 2.490 10.050 2.730 ;
        RECT  6.940 1.130 7.180 3.570 ;
        RECT  5.930 3.330 7.180 3.570 ;
        RECT  2.030 1.740 3.240 1.980 ;
        RECT  3.000 2.600 5.880 2.840 ;
        RECT  5.480 2.600 5.880 3.030 ;
        RECT  2.030 3.240 3.240 3.480 ;
        RECT  3.000 1.740 3.240 3.800 ;
        RECT  9.810 3.380 10.440 3.620 ;
        RECT  3.000 3.560 4.110 3.800 ;
        RECT  9.810 3.360 10.050 4.040 ;
        RECT  9.140 3.800 10.050 4.040 ;
        RECT  3.870 3.560 4.110 4.470 ;
        RECT  9.140 3.800 9.380 4.470 ;
        RECT  3.870 4.230 9.380 4.470 ;
    END
END su01d0

MACRO srlab4
    CLASS CORE ;
    FOREIGN srlab4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.732  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.150 2.010 7.870 2.250 ;
        RECT  7.630 1.570 7.870 2.250 ;
        RECT  7.340 2.010 7.780 2.460 ;
        RECT  7.360 2.010 7.600 4.310 ;
        RECT  6.060 3.720 7.600 3.990 ;
        RECT  6.150 1.560 6.390 2.250 ;
        RECT  6.060 3.720 6.300 4.340 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.531  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.330 2.580 6.100 3.020 ;
        RECT  4.760 3.550 5.570 3.790 ;
        RECT  5.330 1.830 5.570 3.790 ;
        RECT  4.730 1.830 5.570 2.070 ;
        RECT  3.350 4.020 5.000 4.260 ;
        RECT  4.760 3.550 5.000 4.260 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.230 2.440 0.550 2.840 ;
        RECT  0.120 2.580 0.500 3.020 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.460 3.300 2.240 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.840 3.210 8.240 5.600 ;
        RECT  6.730 4.620 7.130 5.600 ;
        RECT  5.420 4.620 5.820 5.600 ;
        RECT  4.110 4.620 4.510 5.600 ;
        RECT  2.800 4.620 3.200 5.600 ;
        RECT  1.460 4.120 1.860 5.600 ;
        RECT  0.150 4.140 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  6.810 0.000 7.210 1.420 ;
        RECT  5.290 0.000 5.690 1.200 ;
        RECT  3.920 0.000 4.320 1.910 ;
        RECT  3.160 0.000 3.560 1.200 ;
        RECT  1.380 0.000 1.780 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.080 0.470 2.200 ;
        RECT  0.230 1.960 1.030 2.200 ;
        RECT  0.790 1.960 1.030 3.560 ;
        RECT  1.710 2.350 2.070 2.750 ;
        RECT  0.790 2.430 1.040 3.560 ;
        RECT  1.710 2.350 1.950 3.130 ;
        RECT  0.790 2.890 1.950 3.130 ;
        RECT  0.790 2.890 1.110 3.560 ;
        RECT  0.720 3.160 1.110 3.560 ;
        RECT  1.270 1.380 2.610 1.620 ;
        RECT  1.270 1.380 1.510 2.010 ;
        RECT  2.370 2.610 5.090 2.850 ;
        RECT  2.370 1.380 2.610 3.760 ;
        RECT  2.030 3.520 2.610 3.760 ;
    END
END srlab4

MACRO srlab2
    CLASS CORE ;
    FOREIGN srlab2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.730  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.020 3.050 6.010 3.450 ;
        RECT  5.670 1.460 6.010 3.450 ;
        RECT  5.100 1.460 6.010 2.170 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.254  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.880 1.460 4.420 2.060 ;
        RECT  3.600 3.050 4.120 3.450 ;
        RECT  3.880 1.460 4.120 3.450 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.050 0.500 3.020 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.610 2.050 2.110 2.450 ;
        RECT  1.820 1.460 2.110 2.450 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.690 4.150 5.930 5.600 ;
        RECT  4.270 4.170 4.510 5.600 ;
        RECT  2.970 4.170 3.210 5.600 ;
        RECT  1.410 4.170 1.650 5.600 ;
        RECT  0.150 4.530 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.770 0.000 5.170 0.980 ;
        RECT  3.080 0.000 3.480 1.220 ;
        RECT  1.430 0.000 1.670 1.150 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.620 2.410 3.630 2.650 ;
        RECT  2.620 1.520 2.870 3.370 ;
        RECT  2.100 3.130 2.870 3.370 ;
        RECT  0.150 1.540 1.060 1.780 ;
        RECT  4.360 2.570 5.270 2.810 ;
        RECT  0.820 1.540 1.060 3.930 ;
        RECT  4.360 2.570 4.600 3.930 ;
        RECT  0.820 3.690 4.600 3.930 ;
        RECT  2.420 3.690 2.660 4.600 ;
    END
END srlab2

MACRO srlab1
    CLASS CORE ;
    FOREIGN srlab1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.240  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.220 1.740 5.280 1.980 ;
        RECT  4.220 1.740 4.460 3.450 ;
        RECT  4.060 2.540 4.460 3.020 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.068  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.520 1.460 3.780 3.450 ;
        RECT  3.400 1.460 3.780 1.960 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.050 0.500 3.020 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.610 2.050 2.110 2.450 ;
        RECT  1.820 1.460 2.110 2.450 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.960 4.170 5.200 5.600 ;
        RECT  2.950 4.190 3.190 5.600 ;
        RECT  1.410 4.170 1.650 5.600 ;
        RECT  0.150 4.530 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.220 0.000 4.460 1.490 ;
        RECT  1.430 0.000 1.670 1.150 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.620 2.090 3.140 2.490 ;
        RECT  2.620 1.520 2.870 3.370 ;
        RECT  2.100 3.130 2.870 3.370 ;
        RECT  0.150 1.540 1.060 1.780 ;
        RECT  0.820 1.540 1.060 3.930 ;
        RECT  4.710 2.520 4.950 3.930 ;
        RECT  0.820 3.690 4.950 3.930 ;
        RECT  2.420 3.690 2.660 4.600 ;
    END
END srlab1

MACRO slnlq4
    CLASS CORE ;
    FOREIGN slnlq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.030 2.050 4.270 2.600 ;
        RECT  3.660 2.360 4.270 2.600 ;
        RECT  3.420 2.580 3.920 3.020 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.860 2.440 17.300 3.020 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.654  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.400 3.060 9.840 3.460 ;
        RECT  9.600 1.910 9.840 3.460 ;
        RECT  7.290 1.910 9.840 2.150 ;
        RECT  8.770 1.240 9.010 2.150 ;
        RECT  8.160 3.060 8.900 3.580 ;
        RECT  7.290 1.240 7.530 2.150 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        RECT  1.970 2.450 2.740 2.690 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.344  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 3.690 16.460 4.120 ;
        RECT  16.200 1.630 16.460 4.120 ;
        RECT  15.850 1.630 16.460 1.870 ;
        RECT  14.840 3.770 16.460 4.010 ;
        RECT  14.840 3.770 15.080 4.350 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.920 5.600 ;
        RECT  16.800 4.310 17.200 5.600 ;
        RECT  15.500 4.620 15.900 5.600 ;
        RECT  14.190 4.620 14.590 5.600 ;
        RECT  12.020 3.890 12.260 5.600 ;
        RECT  9.260 4.390 9.660 5.600 ;
        RECT  7.600 4.350 8.000 5.600 ;
        RECT  6.290 4.400 6.690 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.800 3.550 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.920 0.740 ;
        RECT  16.440 0.000 16.840 0.910 ;
        RECT  15.060 0.000 15.470 0.910 ;
        RECT  12.510 0.000 12.750 1.200 ;
        RECT  9.510 0.000 9.750 1.640 ;
        RECT  8.030 0.000 8.270 1.640 ;
        RECT  6.550 0.000 6.790 1.640 ;
        RECT  3.240 0.000 3.640 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.430 1.250 1.670 ;
        RECT  1.010 1.430 1.250 3.310 ;
        RECT  0.230 3.070 1.250 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.590 1.620 1.830 2.170 ;
        RECT  1.590 1.930 3.390 2.170 ;
        RECT  1.490 1.940 1.730 3.840 ;
        RECT  1.280 3.600 1.520 4.600 ;
        RECT  1.280 4.360 1.860 4.600 ;
        RECT  2.040 1.010 2.710 1.250 ;
        RECT  2.470 1.010 2.710 1.680 ;
        RECT  2.470 1.440 4.790 1.680 ;
        RECT  4.550 1.440 4.790 3.100 ;
        RECT  4.290 2.860 4.790 3.100 ;
        RECT  2.070 3.390 2.810 3.630 ;
        RECT  4.290 2.860 4.530 3.820 ;
        RECT  2.560 3.580 4.530 3.820 ;
        RECT  2.070 3.390 2.310 4.000 ;
        RECT  5.590 1.800 5.830 3.570 ;
        RECT  5.030 0.980 6.310 1.240 ;
        RECT  5.030 0.980 5.490 1.380 ;
        RECT  6.070 0.980 6.310 2.130 ;
        RECT  6.070 1.890 6.920 2.130 ;
        RECT  6.680 1.890 6.920 2.800 ;
        RECT  6.680 2.400 9.360 2.800 ;
        RECT  5.030 0.980 5.270 4.280 ;
        RECT  4.940 3.860 5.360 4.280 ;
        RECT  10.080 1.210 10.580 1.610 ;
        RECT  6.190 2.420 6.430 4.110 ;
        RECT  10.080 1.210 10.320 4.110 ;
        RECT  6.190 3.870 10.320 4.110 ;
        RECT  11.490 0.980 12.090 1.220 ;
        RECT  11.490 0.980 11.730 2.690 ;
        RECT  11.220 2.450 11.730 2.690 ;
        RECT  11.220 2.450 11.460 3.170 ;
        RECT  11.220 2.930 11.770 3.170 ;
        RECT  11.000 1.210 11.240 2.210 ;
        RECT  10.710 1.970 11.240 2.210 ;
        RECT  12.450 1.990 13.030 2.230 ;
        RECT  12.450 1.990 12.690 2.550 ;
        RECT  12.030 2.380 12.650 2.620 ;
        RECT  10.710 1.970 10.950 3.650 ;
        RECT  12.030 2.380 12.270 3.650 ;
        RECT  10.680 3.410 12.270 3.650 ;
        RECT  10.680 3.400 10.920 4.620 ;
        RECT  14.130 1.090 14.370 1.680 ;
        RECT  13.860 1.440 14.370 1.680 ;
        RECT  13.860 1.440 14.100 3.450 ;
        RECT  13.350 3.210 14.100 3.450 ;
        RECT  13.350 3.210 13.810 3.610 ;
        RECT  13.350 3.210 13.590 3.930 ;
        RECT  13.030 3.680 13.450 4.140 ;
        RECT  13.250 1.130 13.490 1.750 ;
        RECT  11.970 1.510 13.610 1.750 ;
        RECT  11.970 1.510 12.210 2.140 ;
        RECT  15.550 2.530 15.960 2.940 ;
        RECT  14.480 2.540 15.960 2.940 ;
        RECT  13.370 1.510 13.610 2.960 ;
        RECT  12.870 2.720 13.610 2.960 ;
        RECT  12.870 2.720 13.110 3.440 ;
        RECT  12.550 3.040 13.110 3.440 ;
        RECT  14.480 2.540 14.720 3.530 ;
        RECT  12.550 3.040 12.790 4.620 ;
        RECT  13.710 4.140 14.580 4.380 ;
        RECT  14.340 3.290 14.580 4.380 ;
        RECT  12.550 4.380 13.950 4.620 ;
        RECT  15.100 1.150 17.800 1.390 ;
        RECT  15.100 1.150 15.340 1.790 ;
        RECT  14.610 1.550 15.340 1.790 ;
        RECT  14.610 1.550 14.850 2.260 ;
        RECT  17.560 1.150 17.800 3.830 ;
        RECT  17.360 3.430 17.800 3.830 ;
    END
END slnlq4

MACRO slnlq2
    CLASS CORE ;
    FOREIGN slnlq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.030 2.050 4.270 2.600 ;
        RECT  3.660 2.360 4.270 2.600 ;
        RECT  3.420 2.580 3.920 3.020 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.620 2.590 15.080 3.030 ;
        RECT  14.630 2.400 15.030 3.030 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.509  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.370 3.060 8.500 3.580 ;
        RECT  8.260 1.830 8.500 3.580 ;
        RECT  7.400 1.830 8.500 2.070 ;
        RECT  7.400 1.550 7.640 2.070 ;
        RECT  7.190 1.240 7.590 1.740 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        RECT  1.970 2.450 2.740 2.690 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.735  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.140 1.850 14.380 2.570 ;
        RECT  13.500 3.140 14.170 3.580 ;
        RECT  13.930 2.330 14.170 3.580 ;
        RECT  13.830 1.850 14.380 2.090 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.680 5.600 ;
        RECT  14.220 4.620 14.620 5.600 ;
        RECT  12.920 4.620 13.320 5.600 ;
        RECT  10.650 3.960 11.050 5.600 ;
        RECT  7.960 4.380 8.360 5.600 ;
        RECT  6.340 4.400 6.760 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.800 3.550 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.680 0.740 ;
        RECT  14.540 0.000 14.940 0.980 ;
        RECT  13.230 0.000 13.630 0.980 ;
        RECT  10.810 0.000 11.210 1.200 ;
        RECT  7.930 1.350 8.550 1.590 ;
        RECT  8.310 0.000 8.550 1.590 ;
        RECT  6.530 0.000 6.770 1.640 ;
        RECT  3.240 0.000 3.640 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.430 1.250 1.670 ;
        RECT  1.010 1.430 1.250 3.310 ;
        RECT  0.230 3.070 1.250 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.590 1.620 1.830 2.170 ;
        RECT  1.590 1.930 3.390 2.170 ;
        RECT  1.490 1.940 1.730 3.840 ;
        RECT  1.280 3.600 1.520 4.600 ;
        RECT  1.280 4.360 1.860 4.600 ;
        RECT  2.040 1.010 2.710 1.250 ;
        RECT  2.470 1.010 2.710 1.690 ;
        RECT  2.470 1.450 4.790 1.690 ;
        RECT  4.550 1.450 4.790 3.100 ;
        RECT  4.290 2.860 4.790 3.100 ;
        RECT  2.070 3.390 2.810 3.630 ;
        RECT  4.290 2.860 4.530 3.820 ;
        RECT  2.560 3.580 4.530 3.820 ;
        RECT  2.070 3.390 2.310 4.000 ;
        RECT  5.570 1.880 5.810 3.240 ;
        RECT  5.590 2.960 5.830 3.570 ;
        RECT  5.090 0.980 5.460 1.390 ;
        RECT  5.090 1.070 6.290 1.310 ;
        RECT  5.090 1.070 5.490 1.390 ;
        RECT  6.050 1.070 6.290 2.220 ;
        RECT  6.050 1.980 6.860 2.220 ;
        RECT  6.620 1.980 6.860 2.550 ;
        RECT  6.620 2.310 8.020 2.550 ;
        RECT  7.070 2.310 8.020 2.730 ;
        RECT  5.090 0.980 5.330 4.280 ;
        RECT  4.940 3.860 5.360 4.280 ;
        RECT  8.790 1.700 9.030 2.340 ;
        RECT  6.140 2.460 6.380 4.140 ;
        RECT  8.810 2.050 9.050 4.140 ;
        RECT  6.140 3.900 9.050 4.140 ;
        RECT  10.120 0.980 10.390 1.530 ;
        RECT  10.120 0.980 10.360 2.380 ;
        RECT  9.930 2.140 10.170 3.130 ;
        RECT  9.930 2.890 10.480 3.130 ;
        RECT  9.300 0.980 9.850 1.220 ;
        RECT  9.610 0.980 9.850 1.700 ;
        RECT  11.080 1.920 11.600 2.240 ;
        RECT  11.080 1.920 11.320 2.620 ;
        RECT  10.770 2.380 11.320 2.620 ;
        RECT  9.440 1.460 9.680 3.030 ;
        RECT  10.770 2.380 11.010 2.900 ;
        RECT  10.720 2.630 10.960 3.610 ;
        RECT  9.390 3.370 10.960 3.610 ;
        RECT  9.390 2.750 9.630 4.620 ;
        RECT  12.330 1.090 12.570 3.580 ;
        RECT  12.150 3.180 12.390 3.830 ;
        RECT  11.860 3.590 12.390 3.830 ;
        RECT  11.860 3.590 12.100 4.140 ;
        RECT  10.630 1.440 12.080 1.680 ;
        RECT  11.630 1.130 11.870 1.680 ;
        RECT  10.600 1.650 10.890 1.770 ;
        RECT  10.600 1.650 10.840 2.140 ;
        RECT  11.670 2.470 12.080 2.710 ;
        RECT  11.840 1.440 12.080 2.710 ;
        RECT  13.290 2.500 13.690 2.900 ;
        RECT  12.990 2.660 13.690 2.900 ;
        RECT  11.560 2.480 11.820 3.250 ;
        RECT  11.420 2.850 11.820 3.250 ;
        RECT  11.370 3.100 11.610 4.620 ;
        RECT  12.420 4.140 13.230 4.380 ;
        RECT  12.990 2.660 13.230 4.380 ;
        RECT  11.370 4.380 12.680 4.620 ;
        RECT  12.810 1.220 15.560 1.460 ;
        RECT  15.130 1.750 15.560 2.150 ;
        RECT  12.810 1.220 13.050 2.270 ;
        RECT  15.320 1.220 15.560 3.540 ;
        RECT  15.000 3.300 15.560 3.540 ;
    END
END slnlq2

MACRO slnlq1
    CLASS CORE ;
    FOREIGN slnlq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.030 1.990 4.270 2.600 ;
        RECT  3.660 2.360 4.270 2.600 ;
        RECT  3.420 2.580 3.920 3.020 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.780 2.580 13.430 3.020 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.168  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.720 2.580 8.410 3.190 ;
        RECT  7.210 3.100 8.360 3.340 ;
        RECT  7.720 2.000 7.960 3.340 ;
        RECT  7.140 1.970 7.840 2.210 ;
        RECT  7.140 1.650 7.540 2.210 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        RECT  1.970 2.450 2.740 2.690 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.370  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.620 2.020 15.000 2.460 ;
        RECT  14.650 1.640 14.890 4.350 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.120 5.600 ;
        RECT  14.000 4.620 14.400 5.600 ;
        RECT  12.810 4.420 13.050 5.600 ;
        RECT  10.490 3.960 10.890 5.600 ;
        RECT  7.800 4.370 8.200 5.600 ;
        RECT  6.340 4.400 6.760 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.800 3.550 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.120 0.740 ;
        RECT  13.980 0.000 14.380 0.980 ;
        RECT  13.290 0.000 13.530 1.090 ;
        RECT  10.920 0.000 11.320 1.200 ;
        RECT  7.960 0.000 8.200 1.760 ;
        RECT  6.590 0.000 6.990 1.260 ;
        RECT  3.240 0.000 3.640 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.430 1.250 1.670 ;
        RECT  1.010 1.430 1.250 3.310 ;
        RECT  0.230 3.070 1.250 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.590 1.620 1.830 2.170 ;
        RECT  1.590 1.930 3.400 2.170 ;
        RECT  1.490 1.940 1.730 3.840 ;
        RECT  1.280 3.600 1.520 4.600 ;
        RECT  1.280 4.360 1.860 4.600 ;
        RECT  2.040 1.010 2.710 1.250 ;
        RECT  2.470 1.010 2.710 1.680 ;
        RECT  4.520 0.980 4.760 1.680 ;
        RECT  2.470 1.440 4.760 1.680 ;
        RECT  4.410 1.440 4.750 1.710 ;
        RECT  4.520 0.980 4.750 3.100 ;
        RECT  4.510 1.440 4.530 3.820 ;
        RECT  4.290 2.860 4.530 3.820 ;
        RECT  2.070 3.390 2.810 3.630 ;
        RECT  2.560 3.580 4.530 3.820 ;
        RECT  2.070 3.390 2.310 4.000 ;
        RECT  5.730 1.710 6.160 2.110 ;
        RECT  5.730 1.710 5.970 2.960 ;
        RECT  5.590 2.720 5.830 3.580 ;
        RECT  5.000 0.990 5.610 1.230 ;
        RECT  6.250 2.450 7.480 2.690 ;
        RECT  5.000 0.990 5.240 4.510 ;
        RECT  6.250 2.450 6.490 4.160 ;
        RECT  5.000 3.920 6.490 4.160 ;
        RECT  5.000 3.920 5.270 4.510 ;
        RECT  8.700 1.650 8.940 3.730 ;
        RECT  6.730 3.070 6.970 4.000 ;
        RECT  8.630 3.290 8.870 4.000 ;
        RECT  6.730 3.760 8.870 4.000 ;
        RECT  10.030 0.980 10.580 1.300 ;
        RECT  10.030 0.980 10.270 1.540 ;
        RECT  9.980 1.380 10.220 2.450 ;
        RECT  10.030 2.290 10.270 3.210 ;
        RECT  9.920 2.810 10.320 3.210 ;
        RECT  9.180 0.980 9.790 1.220 ;
        RECT  10.990 2.050 11.540 2.290 ;
        RECT  10.990 2.050 11.230 2.560 ;
        RECT  10.580 2.380 11.180 2.620 ;
        RECT  9.180 0.980 9.420 3.650 ;
        RECT  10.580 2.380 10.820 3.690 ;
        RECT  9.230 3.450 10.820 3.690 ;
        RECT  9.230 3.450 9.470 4.620 ;
        RECT  12.270 1.090 12.760 1.490 ;
        RECT  11.900 3.180 12.510 3.580 ;
        RECT  12.270 1.090 12.510 3.580 ;
        RECT  11.700 3.490 12.150 3.730 ;
        RECT  11.700 3.490 11.940 4.140 ;
        RECT  12.860 1.720 14.170 1.960 ;
        RECT  13.670 1.720 14.170 2.160 ;
        RECT  12.750 1.730 12.990 2.270 ;
        RECT  13.670 1.720 13.910 3.560 ;
        RECT  13.290 3.320 13.910 3.560 ;
        RECT  10.510 1.570 12.030 1.810 ;
        RECT  11.690 1.130 12.030 1.810 ;
        RECT  10.460 1.690 10.730 2.140 ;
        RECT  11.470 2.610 12.030 2.850 ;
        RECT  11.790 1.130 12.030 2.850 ;
        RECT  11.260 2.850 11.740 2.920 ;
        RECT  11.420 2.770 11.660 3.250 ;
        RECT  11.260 2.850 11.660 3.250 ;
        RECT  13.310 3.840 14.390 4.080 ;
        RECT  14.150 2.530 14.390 4.080 ;
        RECT  12.330 3.940 13.610 4.180 ;
        RECT  11.210 2.980 11.450 4.620 ;
        RECT  12.330 3.940 12.570 4.620 ;
        RECT  11.210 4.380 12.570 4.620 ;
    END
END slnlq1

MACRO slnln4
    CLASS CORE ;
    FOREIGN slnln4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.180 3.020 ;
        RECT  1.760 2.350 2.160 3.020 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.460 3.140 18.920 3.580 ;
        RECT  18.460 2.760 18.860 3.580 ;
        END
    END EN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.819  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.220 1.860 9.080 2.100 ;
        RECT  8.840 1.510 9.080 2.100 ;
        RECT  6.220 3.580 8.770 3.980 ;
        RECT  7.360 1.510 7.600 2.100 ;
        RECT  6.220 3.140 6.660 3.980 ;
        RECT  6.220 1.860 6.570 3.980 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.460 0.540 2.920 ;
        RECT  0.120 2.020 0.500 2.460 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.390 3.020 ;
        RECT  4.150 2.210 4.390 3.020 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.781  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.280 1.440 15.080 1.680 ;
        RECT  14.680 1.070 15.080 1.680 ;
        RECT  12.280 3.220 15.070 3.620 ;
        RECT  13.200 1.070 13.600 1.680 ;
        RECT  12.280 2.580 12.830 3.620 ;
        RECT  12.280 1.440 12.680 3.620 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.040 5.600 ;
        RECT  17.750 4.620 18.150 5.600 ;
        RECT  15.440 4.340 15.840 5.600 ;
        RECT  13.900 4.340 14.300 5.600 ;
        RECT  12.040 4.340 12.440 5.600 ;
        RECT  9.330 4.710 9.730 5.600 ;
        RECT  7.760 4.710 8.160 5.600 ;
        RECT  6.360 4.710 6.760 5.600 ;
        RECT  3.200 4.190 3.600 5.600 ;
        RECT  0.720 4.460 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.040 0.740 ;
        RECT  17.850 0.000 18.250 0.950 ;
        RECT  15.420 0.000 15.820 1.200 ;
        RECT  13.940 0.000 14.340 1.200 ;
        RECT  12.460 0.000 12.860 1.200 ;
        RECT  9.500 0.000 9.900 1.620 ;
        RECT  8.020 0.000 8.420 1.620 ;
        RECT  6.540 0.000 6.940 1.620 ;
        RECT  3.270 0.000 3.670 0.890 ;
        RECT  0.740 0.000 1.140 1.050 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.500 1.020 1.740 ;
        RECT  0.780 2.330 1.480 2.570 ;
        RECT  0.780 1.500 1.020 3.400 ;
        RECT  0.150 3.160 1.020 3.400 ;
        RECT  1.510 1.790 3.180 2.030 ;
        RECT  1.510 1.660 1.910 2.060 ;
        RECT  2.370 3.230 3.180 3.470 ;
        RECT  2.940 1.790 3.180 3.470 ;
        RECT  1.460 3.260 2.600 3.500 ;
        RECT  2.040 0.980 2.620 1.220 ;
        RECT  2.380 0.980 2.620 1.550 ;
        RECT  2.380 1.310 4.870 1.550 ;
        RECT  4.630 1.310 4.870 3.600 ;
        RECT  4.100 3.360 4.870 3.600 ;
        RECT  2.720 3.710 4.340 3.950 ;
        RECT  4.100 3.360 4.340 3.950 ;
        RECT  1.990 3.940 2.960 4.180 ;
        RECT  5.640 1.330 6.200 1.570 ;
        RECT  5.640 1.330 5.880 3.390 ;
        RECT  5.670 3.250 5.910 3.840 ;
        RECT  9.990 2.500 10.230 3.220 ;
        RECT  9.420 2.980 10.230 3.220 ;
        RECT  5.140 1.270 5.380 4.570 ;
        RECT  9.420 2.980 9.660 4.460 ;
        RECT  4.990 4.220 9.660 4.460 ;
        RECT  4.990 4.170 5.390 4.570 ;
        RECT  10.240 1.220 10.710 1.620 ;
        RECT  9.510 2.020 10.710 2.260 ;
        RECT  9.510 2.020 9.750 2.580 ;
        RECT  6.880 2.340 9.750 2.580 ;
        RECT  10.470 1.220 10.710 3.700 ;
        RECT  9.900 3.460 10.710 3.700 ;
        RECT  11.800 1.210 12.040 3.080 ;
        RECT  11.440 2.840 12.040 3.080 ;
        RECT  16.070 0.980 16.780 1.220 ;
        RECT  16.070 0.980 16.310 1.810 ;
        RECT  15.690 1.570 16.310 1.810 ;
        RECT  13.020 1.920 15.930 2.320 ;
        RECT  15.690 1.570 15.930 3.620 ;
        RECT  15.690 3.380 16.410 3.620 ;
        RECT  10.950 1.220 11.380 1.620 ;
        RECT  16.250 2.050 16.490 3.140 ;
        RECT  16.250 2.900 16.890 3.140 ;
        RECT  10.950 3.860 16.890 4.100 ;
        RECT  16.650 2.900 16.890 4.100 ;
        RECT  10.950 1.220 11.190 4.490 ;
        RECT  10.670 4.090 11.190 4.490 ;
        RECT  16.890 2.090 17.400 2.490 ;
        RECT  17.160 1.530 17.400 4.580 ;
        RECT  16.840 4.340 17.400 4.580 ;
        RECT  17.640 1.610 18.840 1.850 ;
        RECT  17.640 1.610 17.890 4.380 ;
        RECT  17.640 4.140 18.890 4.380 ;
    END
END slnln4

MACRO slnln2
    CLASS CORE ;
    FOREIGN slnln2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.180 3.020 ;
        RECT  1.760 2.390 2.160 3.020 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.000 2.020 15.560 2.610 ;
        END
    END EN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.408  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 3.020 7.790 3.260 ;
        RECT  6.780 1.730 7.600 1.970 ;
        RECT  7.360 1.270 7.600 1.970 ;
        RECT  6.780 1.730 7.220 3.260 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.020 0.540 2.920 ;
        RECT  0.120 2.020 0.540 2.460 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.390 3.020 ;
        RECT  4.150 2.210 4.390 3.020 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.444  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.260 2.600 12.120 3.020 ;
        RECT  11.260 1.440 12.040 1.720 ;
        RECT  11.800 1.090 12.040 1.720 ;
        RECT  11.260 1.440 11.700 3.020 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.680 5.600 ;
        RECT  14.390 4.620 14.790 5.600 ;
        RECT  12.510 4.710 12.910 5.600 ;
        RECT  11.150 4.710 11.550 5.600 ;
        RECT  8.040 4.710 8.440 5.600 ;
        RECT  6.620 4.710 7.020 5.600 ;
        RECT  3.190 4.190 3.590 5.600 ;
        RECT  0.720 4.460 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.680 0.740 ;
        RECT  14.540 0.000 14.940 0.950 ;
        RECT  12.540 0.000 12.780 1.220 ;
        RECT  10.980 0.000 11.380 1.200 ;
        RECT  8.020 0.000 8.420 1.510 ;
        RECT  6.540 0.000 6.940 1.490 ;
        RECT  3.270 0.000 3.670 0.890 ;
        RECT  0.740 0.000 1.140 1.050 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.500 1.020 1.740 ;
        RECT  0.780 2.330 1.480 2.570 ;
        RECT  0.780 1.500 1.020 3.400 ;
        RECT  0.150 3.160 1.020 3.400 ;
        RECT  1.510 1.790 3.180 2.030 ;
        RECT  1.510 1.660 1.910 2.060 ;
        RECT  2.370 3.230 3.180 3.470 ;
        RECT  2.940 1.790 3.180 3.470 ;
        RECT  1.460 3.260 2.590 3.500 ;
        RECT  2.040 0.980 2.620 1.220 ;
        RECT  2.380 0.980 2.620 1.550 ;
        RECT  2.380 1.310 4.880 1.550 ;
        RECT  4.640 1.310 4.880 3.600 ;
        RECT  3.990 3.360 4.880 3.600 ;
        RECT  2.710 3.710 4.230 3.950 ;
        RECT  3.990 3.360 4.230 3.950 ;
        RECT  1.990 3.940 2.950 4.180 ;
        RECT  5.800 1.250 6.200 1.650 ;
        RECT  5.960 1.250 6.200 3.350 ;
        RECT  5.960 2.950 6.400 3.350 ;
        RECT  5.140 1.270 5.380 3.940 ;
        RECT  8.400 2.270 8.640 3.940 ;
        RECT  5.140 3.700 8.640 3.940 ;
        RECT  8.840 1.220 9.130 1.990 ;
        RECT  7.840 1.750 9.130 1.990 ;
        RECT  7.840 1.750 8.080 2.610 ;
        RECT  7.640 2.210 8.080 2.610 ;
        RECT  8.890 1.220 9.130 3.430 ;
        RECT  10.320 1.210 10.560 2.510 ;
        RECT  10.350 2.220 10.590 3.190 ;
        RECT  10.350 2.790 10.780 3.190 ;
        RECT  12.880 2.050 13.120 2.840 ;
        RECT  12.480 2.600 13.120 2.840 ;
        RECT  9.580 1.210 9.820 3.760 ;
        RECT  12.480 2.600 12.720 3.760 ;
        RECT  9.580 3.520 12.720 3.760 ;
        RECT  13.040 0.980 13.600 1.220 ;
        RECT  13.040 0.980 13.280 1.810 ;
        RECT  12.300 1.570 13.600 1.810 ;
        RECT  12.300 1.570 12.540 2.360 ;
        RECT  11.970 1.960 12.540 2.360 ;
        RECT  13.360 1.570 13.600 3.490 ;
        RECT  13.080 3.090 13.600 3.490 ;
        RECT  13.850 1.500 14.090 2.480 ;
        RECT  5.840 4.220 14.130 4.460 ;
        RECT  13.890 1.900 14.130 4.460 ;
        RECT  4.770 4.380 6.180 4.620 ;
        RECT  14.520 1.480 15.530 1.720 ;
        RECT  14.370 2.760 14.770 3.160 ;
        RECT  14.520 1.480 14.760 3.650 ;
        RECT  14.520 3.410 15.450 3.650 ;
        RECT  15.210 3.410 15.450 4.570 ;
    END
END slnln2

MACRO slnln1
    CLASS CORE ;
    FOREIGN slnln1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.180 3.020 ;
        RECT  1.760 2.270 2.160 3.020 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.620 2.580 15.260 3.160 ;
        END
    END EN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.169  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.170 2.010 7.600 2.250 ;
        RECT  7.360 1.650 7.600 2.250 ;
        RECT  6.170 3.580 7.360 3.980 ;
        RECT  6.170 2.980 6.660 3.980 ;
        RECT  6.170 2.010 6.410 3.980 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.460 0.540 2.920 ;
        RECT  0.120 2.020 0.500 2.460 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.390 3.020 ;
        RECT  4.150 2.210 4.390 3.020 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.157  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.610 1.490 11.850 1.730 ;
        RECT  11.610 1.140 11.850 1.730 ;
        RECT  10.610 3.370 11.540 3.610 ;
        RECT  10.610 3.140 11.140 3.610 ;
        RECT  10.610 1.490 10.850 3.610 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.680 5.600 ;
        RECT  14.060 4.620 14.460 5.600 ;
        RECT  11.840 4.340 12.240 5.600 ;
        RECT  10.370 4.340 10.770 5.600 ;
        RECT  7.660 4.710 8.060 5.600 ;
        RECT  6.360 4.710 6.760 5.600 ;
        RECT  3.270 4.190 3.510 5.600 ;
        RECT  0.720 4.460 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.680 0.740 ;
        RECT  14.250 0.000 14.650 0.950 ;
        RECT  12.120 0.000 12.520 0.890 ;
        RECT  10.790 0.000 11.190 1.250 ;
        RECT  7.800 0.000 8.200 1.260 ;
        RECT  6.620 0.000 6.860 1.760 ;
        RECT  3.270 0.000 3.670 0.890 ;
        RECT  0.740 0.000 1.140 1.050 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.500 1.020 1.740 ;
        RECT  0.780 2.330 1.480 2.570 ;
        RECT  0.780 1.500 1.020 3.400 ;
        RECT  0.150 3.160 1.020 3.400 ;
        RECT  1.510 1.640 1.910 2.030 ;
        RECT  1.510 1.790 3.180 2.030 ;
        RECT  2.370 3.230 3.180 3.470 ;
        RECT  2.940 1.790 3.180 3.470 ;
        RECT  1.460 3.260 2.590 3.500 ;
        RECT  2.040 0.980 2.620 1.220 ;
        RECT  2.380 1.130 4.640 1.370 ;
        RECT  4.400 1.130 4.640 1.970 ;
        RECT  4.630 1.730 4.870 3.600 ;
        RECT  4.090 3.360 4.870 3.600 ;
        RECT  2.710 3.710 4.330 3.950 ;
        RECT  4.090 3.360 4.330 3.950 ;
        RECT  1.990 3.940 2.950 4.180 ;
        RECT  5.650 1.520 6.200 1.760 ;
        RECT  5.650 1.520 5.890 3.440 ;
        RECT  5.670 3.300 5.910 3.840 ;
        RECT  8.320 2.500 8.560 3.220 ;
        RECT  7.750 2.980 8.560 3.220 ;
        RECT  7.750 2.980 7.990 4.460 ;
        RECT  4.990 4.220 7.990 4.460 ;
        RECT  5.140 1.470 5.380 4.570 ;
        RECT  4.990 4.170 5.380 4.570 ;
        RECT  8.570 1.240 9.040 1.740 ;
        RECT  7.840 1.500 9.040 1.740 ;
        RECT  7.840 1.500 8.080 2.730 ;
        RECT  6.880 2.490 8.080 2.730 ;
        RECT  8.800 1.240 9.040 3.700 ;
        RECT  8.230 3.460 9.040 3.700 ;
        RECT  10.130 1.210 10.370 3.080 ;
        RECT  9.770 2.840 10.370 3.080 ;
        RECT  9.280 1.210 9.710 1.610 ;
        RECT  12.650 2.050 12.890 3.140 ;
        RECT  12.650 2.900 13.290 3.140 ;
        RECT  9.280 3.860 13.290 4.100 ;
        RECT  13.050 2.900 13.290 4.100 ;
        RECT  9.280 1.210 9.520 4.490 ;
        RECT  9.000 4.090 9.520 4.490 ;
        RECT  12.750 0.980 13.310 1.220 ;
        RECT  12.750 0.980 12.990 1.810 ;
        RECT  12.090 1.570 12.990 1.810 ;
        RECT  11.100 1.980 12.330 2.380 ;
        RECT  12.090 1.570 12.330 3.620 ;
        RECT  12.090 3.380 12.810 3.620 ;
        RECT  13.290 2.090 13.800 2.490 ;
        RECT  13.560 1.560 13.800 4.580 ;
        RECT  13.240 4.340 13.800 4.580 ;
        RECT  14.050 1.640 15.240 1.880 ;
        RECT  14.050 1.640 14.290 3.640 ;
        RECT  14.050 3.400 15.210 3.640 ;
    END
END slnln1

MACRO slnlb4
    CLASS CORE ;
    FOREIGN slnlb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.010 2.740 2.460 ;
        RECT  2.410 2.010 2.650 3.060 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 5.190 2.420 ;
        RECT  4.540 2.020 4.980 2.460 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.659  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  20.170 3.130 20.600 3.580 ;
        RECT  20.220 1.570 20.600 3.580 ;
        RECT  19.280 1.570 20.600 1.810 ;
        RECT  18.230 3.130 20.600 3.370 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.260 1.460 18.420 1.900 ;
        RECT  16.250 1.410 18.050 1.650 ;
        RECT  17.650 1.080 18.050 1.900 ;
        RECT  16.390 2.390 17.510 2.630 ;
        RECT  17.260 1.410 17.510 2.630 ;
        RECT  15.590 3.540 17.290 3.780 ;
        RECT  16.390 2.390 16.630 3.780 ;
        RECT  16.250 1.050 16.490 1.650 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.500 0.540 2.830 ;
        RECT  0.120 2.500 0.510 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.980 2.910 1.220 ;
        RECT  1.630 2.660 2.050 3.060 ;
        RECT  1.380 3.140 1.870 3.380 ;
        RECT  1.630 0.980 1.870 3.380 ;
        RECT  1.180 3.700 1.620 4.140 ;
        RECT  1.380 3.140 1.620 4.140 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.180 1.460 15.620 1.900 ;
        RECT  13.570 2.450 15.580 2.690 ;
        RECT  15.340 1.460 15.580 2.690 ;
        RECT  13.290 1.430 15.440 1.670 ;
        RECT  14.770 1.070 15.010 1.670 ;
        RECT  13.290 0.980 13.530 1.670 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.720 5.600 ;
        RECT  20.170 3.900 20.570 5.600 ;
        RECT  18.810 3.810 19.210 5.600 ;
        RECT  17.450 4.610 17.870 5.600 ;
        RECT  16.150 4.610 16.550 5.600 ;
        RECT  14.310 4.610 14.710 5.600 ;
        RECT  13.000 4.610 13.400 5.600 ;
        RECT  11.620 4.710 12.020 5.600 ;
        RECT  8.410 4.380 8.810 5.600 ;
        RECT  5.210 4.290 5.610 5.600 ;
        RECT  3.130 4.490 3.530 5.600 ;
        RECT  0.720 4.530 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.720 0.740 ;
        RECT  20.050 0.000 20.450 1.170 ;
        RECT  18.570 0.000 18.970 1.160 ;
        RECT  16.910 0.000 17.310 0.980 ;
        RECT  15.430 0.000 15.830 0.980 ;
        RECT  13.950 0.000 14.350 0.980 ;
        RECT  11.170 0.000 11.570 0.890 ;
        RECT  9.370 0.000 9.770 0.890 ;
        RECT  5.350 0.000 5.750 0.890 ;
        RECT  3.290 0.000 3.690 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.020 1.820 ;
        RECT  0.780 1.580 1.020 2.420 ;
        RECT  0.780 2.180 1.290 2.420 ;
        RECT  1.050 2.180 1.290 2.900 ;
        RECT  0.780 2.660 1.290 2.900 ;
        RECT  0.780 2.660 1.020 3.520 ;
        RECT  0.150 3.280 1.020 3.520 ;
        RECT  3.460 1.310 4.460 1.550 ;
        RECT  3.460 1.310 3.700 3.520 ;
        RECT  3.460 3.280 4.240 3.520 ;
        RECT  4.760 1.330 5.790 1.570 ;
        RECT  5.550 1.330 5.790 2.920 ;
        RECT  5.470 2.520 5.870 2.920 ;
        RECT  5.290 2.680 5.530 3.370 ;
        RECT  4.540 3.130 5.530 3.370 ;
        RECT  2.110 1.510 3.220 1.750 ;
        RECT  2.980 1.510 3.220 4.000 ;
        RECT  6.060 3.660 7.140 3.900 ;
        RECT  6.900 1.460 7.140 3.900 ;
        RECT  1.920 3.760 6.300 4.000 ;
        RECT  8.200 1.460 8.700 1.780 ;
        RECT  8.200 1.460 8.440 2.260 ;
        RECT  7.860 2.020 8.440 2.260 ;
        RECT  7.860 2.020 8.100 3.450 ;
        RECT  7.860 3.050 8.280 3.450 ;
        RECT  6.200 1.050 9.190 1.220 ;
        RECT  6.200 0.980 9.130 1.220 ;
        RECT  8.890 1.130 10.420 1.290 ;
        RECT  8.950 1.130 10.420 1.370 ;
        RECT  6.200 0.980 6.440 2.310 ;
        RECT  6.260 2.150 6.500 3.400 ;
        RECT  5.840 3.160 6.500 3.400 ;
        RECT  11.140 1.610 11.540 1.930 ;
        RECT  11.140 1.610 11.380 3.510 ;
        RECT  10.980 3.110 11.380 3.510 ;
        RECT  10.660 1.130 12.050 1.370 ;
        RECT  11.810 1.130 12.050 1.930 ;
        RECT  10.660 1.130 10.900 1.790 ;
        RECT  11.810 1.690 12.340 1.930 ;
        RECT  10.400 1.620 10.820 2.020 ;
        RECT  12.100 1.690 12.340 2.290 ;
        RECT  12.320 2.050 12.560 2.610 ;
        RECT  10.580 1.550 10.820 2.900 ;
        RECT  10.320 2.660 10.820 2.900 ;
        RECT  10.320 2.660 10.560 3.500 ;
        RECT  12.590 0.980 12.830 1.810 ;
        RECT  12.800 1.910 14.570 2.150 ;
        RECT  11.620 2.170 11.860 3.370 ;
        RECT  12.800 1.570 13.040 3.370 ;
        RECT  11.620 3.130 13.040 3.370 ;
        RECT  8.940 1.660 10.080 2.060 ;
        RECT  15.900 1.900 17.020 2.150 ;
        RECT  8.680 2.020 9.180 2.260 ;
        RECT  8.680 2.020 8.920 2.740 ;
        RECT  8.340 2.500 8.920 2.740 ;
        RECT  15.900 1.900 16.140 3.170 ;
        RECT  13.310 2.930 16.140 3.170 ;
        RECT  9.490 3.480 10.080 3.720 ;
        RECT  9.840 1.660 10.080 3.990 ;
        RECT  11.620 3.610 13.550 3.850 ;
        RECT  13.310 2.930 13.550 3.850 ;
        RECT  9.840 3.750 11.860 3.990 ;
        RECT  7.380 1.540 7.960 1.780 ;
        RECT  17.750 2.520 19.800 2.760 ;
        RECT  9.160 2.520 9.400 3.220 ;
        RECT  8.520 2.980 9.400 3.220 ;
        RECT  7.380 1.540 7.620 3.930 ;
        RECT  8.520 2.980 8.760 4.140 ;
        RECT  7.380 3.690 7.980 3.930 ;
        RECT  7.740 3.900 9.330 4.140 ;
        RECT  12.070 4.120 17.990 4.360 ;
        RECT  17.750 2.520 17.990 4.360 ;
        RECT  9.090 3.900 9.330 4.620 ;
        RECT  10.710 4.230 12.310 4.470 ;
        RECT  7.740 3.690 7.980 4.620 ;
        RECT  7.100 4.380 7.980 4.620 ;
        RECT  9.090 4.380 10.950 4.620 ;
    END
END slnlb4

MACRO slnlb2
    CLASS CORE ;
    FOREIGN slnlb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.010 2.740 2.460 ;
        RECT  2.430 2.010 2.670 3.060 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 5.090 2.460 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.493  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.270 1.460 16.740 1.900 ;
        RECT  16.270 1.460 16.510 4.300 ;
        RECT  15.840 1.460 16.740 1.700 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.530  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.890 3.570 15.360 3.890 ;
        RECT  15.120 1.380 15.360 3.890 ;
        RECT  14.620 1.380 15.360 1.900 ;
        RECT  14.510 1.380 15.360 1.700 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.500 0.540 2.830 ;
        RECT  0.120 2.500 0.510 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.980 2.930 1.220 ;
        RECT  1.630 2.660 2.070 3.060 ;
        RECT  1.380 3.140 1.870 3.380 ;
        RECT  1.630 0.980 1.870 3.380 ;
        RECT  1.180 3.700 1.620 4.140 ;
        RECT  1.380 3.140 1.620 4.140 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.646  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.670 1.730 14.210 2.130 ;
        RECT  13.500 1.460 13.940 1.900 ;
        RECT  13.670 1.460 13.910 3.410 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.360 5.600 ;
        RECT  16.870 3.130 17.110 5.600 ;
        RECT  15.630 4.610 16.030 5.600 ;
        RECT  14.330 4.610 14.730 5.600 ;
        RECT  13.020 4.610 13.420 5.600 ;
        RECT  11.720 4.710 12.120 5.600 ;
        RECT  8.410 4.380 8.810 5.600 ;
        RECT  5.210 4.290 5.610 5.600 ;
        RECT  3.130 4.490 3.530 5.600 ;
        RECT  0.720 4.530 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.360 0.740 ;
        RECT  15.250 0.000 15.650 0.980 ;
        RECT  13.030 0.000 13.430 0.890 ;
        RECT  12.330 0.000 12.730 0.890 ;
        RECT  9.370 0.000 9.770 0.890 ;
        RECT  5.370 0.000 5.770 0.890 ;
        RECT  3.310 0.000 3.710 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.020 1.820 ;
        RECT  0.780 1.580 1.020 2.420 ;
        RECT  0.780 2.180 1.310 2.420 ;
        RECT  1.070 2.180 1.310 2.900 ;
        RECT  0.780 2.660 1.310 2.900 ;
        RECT  0.780 2.660 1.020 3.520 ;
        RECT  0.150 3.280 1.020 3.520 ;
        RECT  3.460 1.310 4.480 1.550 ;
        RECT  3.460 1.310 3.700 3.520 ;
        RECT  3.460 3.280 4.240 3.520 ;
        RECT  4.780 1.330 5.790 1.570 ;
        RECT  5.550 1.330 5.790 2.920 ;
        RECT  5.470 2.520 5.870 2.920 ;
        RECT  5.290 2.600 5.530 3.370 ;
        RECT  4.540 3.130 5.530 3.370 ;
        RECT  2.110 1.510 3.220 1.750 ;
        RECT  2.980 1.510 3.220 4.000 ;
        RECT  6.060 3.660 7.160 3.900 ;
        RECT  6.920 1.460 7.160 3.900 ;
        RECT  1.920 3.760 6.300 4.000 ;
        RECT  8.220 1.460 8.720 1.780 ;
        RECT  8.220 1.460 8.460 2.260 ;
        RECT  7.880 2.020 8.460 2.260 ;
        RECT  7.880 2.020 8.120 3.450 ;
        RECT  7.880 3.050 8.280 3.450 ;
        RECT  6.220 1.050 9.190 1.220 ;
        RECT  6.220 0.980 9.130 1.220 ;
        RECT  8.890 1.130 10.440 1.290 ;
        RECT  8.950 1.130 10.440 1.370 ;
        RECT  6.220 0.980 6.460 2.380 ;
        RECT  6.250 2.260 6.490 3.400 ;
        RECT  5.840 3.160 6.490 3.400 ;
        RECT  11.160 1.600 11.560 1.920 ;
        RECT  11.160 1.600 11.400 3.510 ;
        RECT  11.020 3.110 11.400 3.510 ;
        RECT  10.680 1.100 12.050 1.340 ;
        RECT  11.810 1.100 12.050 1.930 ;
        RECT  11.810 1.690 12.340 1.930 ;
        RECT  10.420 1.620 10.920 2.020 ;
        RECT  12.100 1.830 12.560 2.070 ;
        RECT  12.320 1.830 12.560 2.610 ;
        RECT  10.680 1.100 10.920 2.890 ;
        RECT  10.330 2.650 10.920 2.890 ;
        RECT  10.330 2.650 10.570 3.500 ;
        RECT  12.540 1.230 13.040 1.550 ;
        RECT  12.800 2.420 13.430 2.820 ;
        RECT  11.640 2.170 11.880 3.370 ;
        RECT  12.800 1.230 13.040 3.370 ;
        RECT  11.640 3.130 13.040 3.370 ;
        RECT  8.960 1.660 10.090 1.980 ;
        RECT  8.960 1.660 9.200 2.260 ;
        RECT  8.700 2.020 9.200 2.260 ;
        RECT  8.700 2.020 8.940 2.740 ;
        RECT  8.360 2.500 8.940 2.740 ;
        RECT  14.640 2.480 14.880 3.330 ;
        RECT  9.510 3.450 10.090 3.690 ;
        RECT  9.850 1.660 10.090 3.990 ;
        RECT  14.410 3.090 14.650 3.890 ;
        RECT  11.600 3.650 14.650 3.890 ;
        RECT  9.850 3.750 11.840 3.990 ;
        RECT  7.400 1.460 7.980 1.780 ;
        RECT  9.180 2.520 9.420 3.220 ;
        RECT  8.520 2.980 9.420 3.220 ;
        RECT  7.400 1.460 7.640 4.140 ;
        RECT  8.520 2.980 8.760 4.140 ;
        RECT  7.400 3.900 9.390 4.140 ;
        RECT  9.150 3.900 9.390 4.470 ;
        RECT  12.060 4.130 15.840 4.370 ;
        RECT  15.600 2.010 15.840 4.370 ;
        RECT  9.150 4.230 12.300 4.470 ;
        RECT  7.440 3.900 7.680 4.620 ;
        RECT  7.100 4.380 7.680 4.620 ;
    END
END slnlb2

MACRO slnlb1
    CLASS CORE ;
    FOREIGN slnlb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.010 2.740 2.460 ;
        RECT  2.430 2.010 2.670 3.060 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 5.170 2.460 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.184  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.680 3.800 16.120 4.120 ;
        RECT  15.880 1.830 16.120 4.120 ;
        RECT  15.740 2.580 16.120 3.020 ;
        RECT  15.330 1.830 16.120 2.070 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.510 1.460 15.060 1.900 ;
        RECT  14.400 1.230 14.800 1.630 ;
        RECT  14.510 1.230 14.750 3.020 ;
        RECT  14.440 2.850 14.680 3.710 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.500 0.540 2.830 ;
        RECT  0.120 2.500 0.510 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.980 2.930 1.220 ;
        RECT  1.630 2.660 2.070 3.060 ;
        RECT  1.380 3.140 1.870 3.380 ;
        RECT  1.630 0.980 1.870 3.380 ;
        RECT  1.180 3.700 1.620 4.140 ;
        RECT  1.380 3.140 1.620 4.140 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.139  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.380 1.460 13.940 1.900 ;
        RECT  13.060 3.270 13.620 3.510 ;
        RECT  13.380 1.020 13.620 3.510 ;
        RECT  13.050 1.020 13.620 1.260 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  15.060 4.710 15.460 5.600 ;
        RECT  13.660 4.710 14.060 5.600 ;
        RECT  11.660 4.710 12.060 5.600 ;
        RECT  8.430 4.380 8.830 5.600 ;
        RECT  5.210 4.290 5.610 5.600 ;
        RECT  3.130 4.490 3.530 5.600 ;
        RECT  0.720 4.530 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  15.330 0.000 15.730 1.150 ;
        RECT  13.830 0.000 14.230 0.890 ;
        RECT  11.930 0.000 12.330 0.890 ;
        RECT  9.420 0.000 9.820 0.890 ;
        RECT  5.370 0.000 5.770 0.890 ;
        RECT  3.310 0.000 3.710 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.020 1.820 ;
        RECT  0.780 1.580 1.020 2.420 ;
        RECT  0.980 2.180 1.310 2.900 ;
        RECT  0.780 2.660 1.020 3.520 ;
        RECT  0.150 3.280 1.020 3.520 ;
        RECT  3.460 1.310 4.480 1.550 ;
        RECT  3.460 1.310 3.700 3.520 ;
        RECT  3.460 3.280 4.240 3.520 ;
        RECT  4.780 1.330 5.790 1.570 ;
        RECT  5.550 1.330 5.790 2.920 ;
        RECT  5.470 2.520 5.870 2.920 ;
        RECT  5.290 2.670 5.530 3.520 ;
        RECT  4.540 3.280 5.530 3.520 ;
        RECT  2.110 1.510 3.220 1.750 ;
        RECT  2.980 1.510 3.220 4.000 ;
        RECT  6.060 3.660 7.160 3.900 ;
        RECT  6.920 1.460 7.160 3.900 ;
        RECT  1.920 3.760 6.300 4.000 ;
        RECT  8.220 1.460 8.720 1.800 ;
        RECT  8.220 1.460 8.460 2.260 ;
        RECT  7.880 2.020 8.460 2.260 ;
        RECT  7.880 2.020 8.120 3.460 ;
        RECT  7.880 3.140 8.320 3.460 ;
        RECT  6.220 0.980 9.190 1.220 ;
        RECT  8.950 1.130 10.440 1.370 ;
        RECT  6.220 0.980 6.460 2.190 ;
        RECT  6.260 2.040 6.500 3.400 ;
        RECT  5.840 3.160 6.500 3.400 ;
        RECT  11.160 1.620 11.560 1.940 ;
        RECT  11.160 1.620 11.400 2.500 ;
        RECT  11.110 2.260 11.350 3.500 ;
        RECT  10.680 1.130 12.360 1.370 ;
        RECT  10.680 1.130 10.920 2.020 ;
        RECT  10.370 1.620 10.920 2.020 ;
        RECT  12.120 1.130 12.360 2.570 ;
        RECT  12.120 2.250 12.640 2.570 ;
        RECT  10.370 1.620 10.610 3.500 ;
        RECT  12.600 1.640 13.120 1.960 ;
        RECT  11.640 2.210 11.880 3.050 ;
        RECT  12.760 2.790 13.120 3.030 ;
        RECT  12.880 1.640 13.120 3.030 ;
        RECT  11.640 2.810 12.960 3.050 ;
        RECT  12.440 2.810 12.680 3.510 ;
        RECT  8.990 1.650 10.130 1.980 ;
        RECT  8.990 1.650 9.230 2.280 ;
        RECT  8.730 2.040 9.230 2.280 ;
        RECT  13.900 2.140 14.270 2.540 ;
        RECT  8.730 2.040 8.970 2.750 ;
        RECT  8.360 2.510 8.970 2.750 ;
        RECT  9.550 3.470 10.130 3.710 ;
        RECT  9.890 1.650 10.130 3.990 ;
        RECT  13.900 2.140 14.150 3.990 ;
        RECT  9.890 3.750 14.150 3.990 ;
        RECT  7.400 1.460 7.980 1.780 ;
        RECT  9.230 2.520 9.470 3.230 ;
        RECT  8.600 2.990 9.470 3.230 ;
        RECT  15.070 2.530 15.310 3.500 ;
        RECT  8.600 2.990 8.840 4.140 ;
        RECT  7.400 1.460 7.640 4.110 ;
        RECT  7.450 3.900 9.380 4.140 ;
        RECT  9.140 3.900 9.380 4.470 ;
        RECT  14.930 3.260 15.170 4.470 ;
        RECT  9.140 4.230 15.170 4.470 ;
        RECT  7.450 3.900 7.690 4.620 ;
        RECT  7.100 4.380 7.690 4.620 ;
    END
END slnlb1

MACRO slnht4
    CLASS CORE ;
    FOREIGN slnht4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.453  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.420 2.580 10.020 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  22.460 2.180 22.840 3.020 ;
        RECT  22.130 2.180 22.840 2.580 ;
        END
    END E
    PIN OE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.499  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.960 1.060 2.460 ;
        END
    END OE
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.210 2.450 7.700 3.080 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.640 2.580 11.230 3.020 ;
        RECT  10.990 2.220 11.230 3.020 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.023  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.730 1.450 19.290 1.690 ;
        RECT  19.050 1.060 19.290 1.690 ;
        RECT  16.730 3.010 18.940 3.410 ;
        RECT  17.570 1.070 17.810 1.690 ;
        RECT  16.730 2.580 17.330 3.410 ;
        RECT  16.730 1.450 16.970 3.410 ;
        END
    END SO
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.987  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.570 1.440 3.430 1.680 ;
        RECT  3.190 0.980 3.430 1.680 ;
        RECT  1.480 3.100 3.190 3.500 ;
        RECT  1.570 1.440 2.180 2.470 ;
        RECT  1.570 1.300 2.030 2.470 ;
        RECT  1.570 1.300 1.810 3.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 22.960 5.600 ;
        RECT  21.630 4.310 21.870 5.600 ;
        RECT  19.140 4.710 19.540 5.600 ;
        RECT  17.770 4.710 18.170 5.600 ;
        RECT  16.300 4.710 16.700 5.600 ;
        RECT  14.870 4.740 15.270 5.600 ;
        RECT  13.520 4.245 13.860 5.600 ;
        RECT  10.270 4.520 10.670 5.600 ;
        RECT  7.790 4.620 8.190 5.600 ;
        RECT  4.710 4.420 4.950 5.600 ;
        RECT  3.350 4.620 3.750 5.600 ;
        RECT  2.050 4.620 2.450 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 22.960 0.740 ;
        RECT  21.750 0.000 21.990 1.440 ;
        RECT  19.950 0.000 20.350 0.890 ;
        RECT  18.310 0.000 18.550 1.200 ;
        RECT  16.830 0.000 17.070 1.210 ;
        RECT  13.645 0.000 14.045 0.840 ;
        RECT  10.190 0.000 10.430 1.310 ;
        RECT  7.670 0.000 8.070 0.890 ;
        RECT  5.580 0.000 5.980 0.890 ;
        RECT  2.450 0.000 2.690 1.200 ;
        RECT  0.970 0.000 1.210 1.200 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.070 0.550 1.470 ;
        RECT  4.630 2.410 5.960 2.650 ;
        RECT  0.120 1.070 0.360 4.000 ;
        RECT  0.120 3.060 0.560 4.000 ;
        RECT  4.630 2.410 4.870 4.000 ;
        RECT  0.120 3.760 4.870 4.000 ;
        RECT  4.150 1.930 6.440 2.170 ;
        RECT  3.300 2.580 4.390 2.820 ;
        RECT  6.200 1.930 6.440 3.180 ;
        RECT  5.370 2.940 6.440 3.180 ;
        RECT  4.150 1.460 4.390 3.260 ;
        RECT  4.140 2.580 4.390 3.260 ;
        RECT  3.670 0.980 5.140 1.220 ;
        RECT  6.380 1.040 6.920 1.570 ;
        RECT  4.810 1.130 6.920 1.570 ;
        RECT  3.670 0.980 3.910 2.160 ;
        RECT  2.610 1.920 3.910 2.160 ;
        RECT  6.680 1.040 6.920 3.760 ;
        RECT  6.060 3.520 6.920 3.760 ;
        RECT  7.160 1.230 7.400 1.820 ;
        RECT  7.160 1.580 8.180 1.820 ;
        RECT  7.940 2.340 8.440 2.740 ;
        RECT  7.940 1.580 8.180 3.590 ;
        RECT  7.160 3.350 8.180 3.590 ;
        RECT  8.440 1.840 9.000 2.080 ;
        RECT  8.760 2.100 10.520 2.340 ;
        RECT  8.760 1.840 9.000 3.140 ;
        RECT  8.620 2.900 8.860 3.670 ;
        RECT  8.460 3.270 8.860 3.670 ;
        RECT  8.910 0.980 9.940 1.220 ;
        RECT  9.700 0.980 9.940 1.790 ;
        RECT  11.310 1.140 11.720 1.790 ;
        RECT  9.700 1.550 11.720 1.790 ;
        RECT  11.470 1.140 11.720 3.600 ;
        RECT  11.400 3.200 11.800 3.600 ;
        RECT  9.160 3.360 11.800 3.600 ;
        RECT  9.160 3.360 9.560 3.760 ;
        RECT  12.850 1.540 13.190 1.845 ;
        RECT  12.900 1.540 13.140 3.075 ;
        RECT  12.900 2.790 13.260 3.075 ;
        RECT  12.040 1.070 14.200 1.310 ;
        RECT  12.040 1.070 12.470 1.560 ;
        RECT  13.960 1.070 14.200 2.450 ;
        RECT  13.960 2.030 14.320 2.450 ;
        RECT  12.230 1.070 12.470 3.075 ;
        RECT  12.180 2.790 12.520 3.075 ;
        RECT  13.370 2.030 13.730 2.450 ;
        RECT  13.490 2.030 13.730 3.545 ;
        RECT  14.550 1.310 14.790 3.545 ;
        RECT  12.235 3.305 14.790 3.545 ;
        RECT  9.790 3.900 12.475 4.140 ;
        RECT  12.235 3.305 12.475 4.140 ;
        RECT  7.290 4.130 10.030 4.370 ;
        RECT  7.290 4.130 7.530 4.620 ;
        RECT  6.330 4.380 7.530 4.620 ;
        RECT  16.090 0.980 16.330 3.500 ;
        RECT  15.740 3.230 16.330 3.500 ;
        RECT  19.620 1.310 20.440 1.550 ;
        RECT  19.620 1.310 19.860 2.260 ;
        RECT  17.660 1.940 19.720 2.340 ;
        RECT  19.480 1.940 19.720 3.260 ;
        RECT  19.480 3.020 20.310 3.260 ;
        RECT  19.960 2.490 20.790 2.730 ;
        RECT  15.350 1.010 15.590 2.990 ;
        RECT  15.050 2.750 15.590 2.990 ;
        RECT  15.050 2.750 15.290 3.980 ;
        RECT  20.550 2.490 20.790 3.980 ;
        RECT  15.050 3.740 20.790 3.980 ;
        RECT  20.920 1.030 21.340 1.440 ;
        RECT  12.960 3.775 14.770 4.015 ;
        RECT  14.530 3.775 14.770 4.470 ;
        RECT  21.030 1.030 21.270 4.470 ;
        RECT  14.530 4.230 21.270 4.470 ;
        RECT  12.960 3.775 13.200 4.620 ;
        RECT  12.380 4.380 13.200 4.620 ;
        RECT  22.490 1.260 22.730 1.920 ;
        RECT  21.530 1.680 22.730 1.920 ;
        RECT  21.530 1.680 21.770 3.510 ;
        RECT  21.530 3.270 22.680 3.510 ;
    END
END slnht4

MACRO slnht2
    CLASS CORE ;
    FOREIGN slnht2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.453  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.120 2.580 8.900 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.650 2.180 20.100 3.020 ;
        END
    END E
    PIN OE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.499  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.630 1.060 2.460 ;
        END
    END OE
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.340 2.140 7.220 2.460 ;
        RECT  6.700 2.020 7.220 2.460 ;
        RECT  6.340 2.140 6.580 2.770 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.340 2.580 10.020 3.020 ;
        RECT  9.610 2.210 10.020 3.020 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.515  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.430 1.450 16.590 1.690 ;
        RECT  16.350 1.070 16.590 1.690 ;
        RECT  15.180 3.090 16.270 3.350 ;
        RECT  15.180 2.570 15.670 3.350 ;
        RECT  15.430 1.450 15.670 3.350 ;
        END
    END SO
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.570  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.710 0.980 1.950 1.520 ;
        RECT  1.180 3.100 1.890 3.590 ;
        RECT  1.550 1.290 1.790 3.590 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.720 5.600 ;
        RECT  18.880 4.300 19.280 5.600 ;
        RECT  16.470 4.710 16.870 5.600 ;
        RECT  15.000 4.710 15.400 5.600 ;
        RECT  13.570 4.740 13.970 5.600 ;
        RECT  12.190 4.360 12.590 5.600 ;
        RECT  8.970 4.520 9.370 5.600 ;
        RECT  6.490 4.620 6.890 5.600 ;
        RECT  3.330 4.420 3.730 5.600 ;
        RECT  2.050 4.620 2.450 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.720 0.740 ;
        RECT  19.190 0.000 19.590 1.440 ;
        RECT  17.010 0.000 17.410 1.200 ;
        RECT  15.530 0.000 15.930 1.210 ;
        RECT  12.335 0.000 12.910 0.820 ;
        RECT  8.890 0.000 9.290 1.310 ;
        RECT  4.100 0.000 4.500 0.890 ;
        RECT  0.890 0.000 1.290 1.200 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 0.980 0.550 1.390 ;
        RECT  3.320 2.410 4.660 2.650 ;
        RECT  0.120 0.980 0.360 3.490 ;
        RECT  0.120 3.060 0.560 3.490 ;
        RECT  0.230 3.060 0.470 4.160 ;
        RECT  3.320 2.410 3.560 4.160 ;
        RECT  0.230 3.920 3.560 4.160 ;
        RECT  2.670 1.930 5.140 2.170 ;
        RECT  2.420 2.440 2.910 2.840 ;
        RECT  2.670 1.460 2.910 2.840 ;
        RECT  4.900 1.930 5.140 3.290 ;
        RECT  4.070 3.050 5.140 3.290 ;
        RECT  2.840 2.500 3.080 3.370 ;
        RECT  2.190 0.980 3.660 1.220 ;
        RECT  3.330 1.130 5.620 1.370 ;
        RECT  3.330 1.130 3.730 1.570 ;
        RECT  2.190 0.980 2.430 2.160 ;
        RECT  2.030 1.760 2.430 2.160 ;
        RECT  5.380 1.130 5.620 3.970 ;
        RECT  4.760 3.730 5.620 3.970 ;
        RECT  5.940 0.980 7.380 1.220 ;
        RECT  5.940 0.980 6.180 1.900 ;
        RECT  5.860 1.490 6.270 1.900 ;
        RECT  5.860 1.490 6.100 3.680 ;
        RECT  5.860 3.270 6.270 3.680 ;
        RECT  7.460 2.100 9.220 2.340 ;
        RECT  7.460 1.770 7.700 3.070 ;
        RECT  7.240 2.830 7.480 3.670 ;
        RECT  7.690 0.980 8.480 1.220 ;
        RECT  8.240 0.980 8.480 1.790 ;
        RECT  10.170 1.140 10.410 1.790 ;
        RECT  8.240 1.550 10.525 1.790 ;
        RECT  10.280 1.550 10.525 3.570 ;
        RECT  7.860 3.330 10.525 3.570 ;
        RECT  11.660 1.540 11.920 3.160 ;
        RECT  10.910 1.060 12.960 1.300 ;
        RECT  12.730 1.060 12.960 2.520 ;
        RECT  12.730 2.100 13.110 2.520 ;
        RECT  10.910 1.060 11.170 3.160 ;
        RECT  13.330 1.230 13.590 1.775 ;
        RECT  13.350 1.230 13.590 3.035 ;
        RECT  12.150 2.160 12.390 3.640 ;
        RECT  13.270 2.795 13.510 3.640 ;
        RECT  10.860 3.400 13.510 3.640 ;
        RECT  7.730 3.810 11.100 4.050 ;
        RECT  10.860 3.400 11.100 4.050 ;
        RECT  5.890 4.000 7.970 4.240 ;
        RECT  5.890 4.000 6.130 4.620 ;
        RECT  5.030 4.380 6.130 4.620 ;
        RECT  14.870 0.980 15.110 2.110 ;
        RECT  14.700 1.830 14.940 3.510 ;
        RECT  14.490 3.110 14.940 3.510 ;
        RECT  17.830 1.070 18.070 1.680 ;
        RECT  16.830 1.440 18.070 1.680 ;
        RECT  16.830 1.440 17.070 2.180 ;
        RECT  16.150 1.940 17.070 2.180 ;
        RECT  16.150 1.940 16.550 2.340 ;
        RECT  16.230 1.940 16.550 2.770 ;
        RECT  16.230 2.530 17.070 2.770 ;
        RECT  16.830 2.530 17.070 3.170 ;
        RECT  16.830 2.930 17.640 3.170 ;
        RECT  14.020 0.980 14.370 1.390 ;
        RECT  17.380 2.140 18.120 2.380 ;
        RECT  14.020 0.980 14.260 3.990 ;
        RECT  13.750 3.340 14.260 3.990 ;
        RECT  17.880 2.140 18.120 3.990 ;
        RECT  13.750 3.750 18.120 3.990 ;
        RECT  18.530 1.030 18.770 3.710 ;
        RECT  11.510 3.880 13.490 4.120 ;
        RECT  13.250 3.880 13.490 4.470 ;
        RECT  18.360 3.460 18.610 4.470 ;
        RECT  13.250 4.230 18.610 4.470 ;
        RECT  11.510 3.880 11.750 4.620 ;
        RECT  11.090 4.380 11.750 4.620 ;
        RECT  20.010 1.240 20.250 1.920 ;
        RECT  19.050 1.680 20.250 1.920 ;
        RECT  19.050 1.680 19.290 3.510 ;
        RECT  19.050 3.270 20.010 3.510 ;
    END
END slnht2

MACRO slnht1
    CLASS CORE ;
    FOREIGN slnht1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.453  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.010 2.580 6.660 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.820 2.180 18.360 3.020 ;
        RECT  17.630 2.180 18.360 2.610 ;
        END
    END E
    PIN OE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.499  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.960 1.060 2.460 ;
        RECT  0.600 1.720 0.960 2.460 ;
        END
    END OE
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.890 2.580 4.460 3.070 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.580 7.930 3.020 ;
        RECT  7.680 2.210 7.930 3.020 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.129  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.290 1.530 16.180 1.920 ;
        RECT  15.740 1.070 16.180 1.920 ;
        RECT  14.980 2.850 15.530 3.170 ;
        RECT  15.290 1.530 15.530 3.170 ;
        END
    END SO
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.529  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.950 2.730 2.830 2.970 ;
        RECT  2.590 1.070 2.830 2.970 ;
        RECT  2.090 1.070 2.830 1.960 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 18.480 5.600 ;
        RECT  16.250 4.300 16.650 5.600 ;
        RECT  14.410 4.400 14.810 5.600 ;
        RECT  13.000 4.710 13.400 5.600 ;
        RECT  11.460 4.750 12.070 5.600 ;
        RECT  10.190 4.240 10.590 5.600 ;
        RECT  6.970 4.520 7.370 5.600 ;
        RECT  4.490 4.620 4.890 5.600 ;
        RECT  3.150 4.270 3.550 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 18.480 0.740 ;
        RECT  17.150 0.000 17.550 1.440 ;
        RECT  14.970 0.000 15.370 1.200 ;
        RECT  13.530 0.000 13.930 1.210 ;
        RECT  11.040 0.000 11.440 0.890 ;
        RECT  6.890 0.000 7.290 1.310 ;
        RECT  4.450 0.000 4.850 0.890 ;
        RECT  3.320 0.000 3.720 0.890 ;
        RECT  0.890 0.000 1.290 1.200 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.060 0.550 1.470 ;
        RECT  1.470 2.200 2.350 2.440 ;
        RECT  0.120 1.060 0.360 3.490 ;
        RECT  1.470 2.200 1.710 3.410 ;
        RECT  0.120 3.170 1.710 3.410 ;
        RECT  0.120 3.090 0.550 3.490 ;
        RECT  3.940 1.230 4.180 1.820 ;
        RECT  3.940 1.580 5.050 1.820 ;
        RECT  4.810 1.580 5.050 2.910 ;
        RECT  4.710 2.700 4.950 3.550 ;
        RECT  3.860 3.310 4.950 3.550 ;
        RECT  5.300 2.100 7.220 2.340 ;
        RECT  5.300 1.760 5.540 3.230 ;
        RECT  5.240 3.070 5.480 3.670 ;
        RECT  5.690 0.980 6.480 1.220 ;
        RECT  6.240 0.980 6.480 1.790 ;
        RECT  6.240 1.550 8.410 1.790 ;
        RECT  8.170 1.140 8.410 3.570 ;
        RECT  8.170 3.170 8.500 3.570 ;
        RECT  5.860 3.330 8.500 3.570 ;
        RECT  9.660 1.510 9.920 3.510 ;
        RECT  10.160 1.680 11.410 1.920 ;
        RECT  10.160 1.680 10.400 3.420 ;
        RECT  10.160 3.180 11.330 3.420 ;
        RECT  8.910 0.990 10.490 1.230 ;
        RECT  10.240 1.150 11.890 1.390 ;
        RECT  11.650 1.150 11.890 2.500 ;
        RECT  10.750 2.250 11.890 2.500 ;
        RECT  3.070 2.120 3.310 4.030 ;
        RECT  5.730 3.810 9.170 4.050 ;
        RECT  3.070 3.790 4.260 4.030 ;
        RECT  8.910 0.990 9.170 4.050 ;
        RECT  4.020 3.910 5.970 4.150 ;
        RECT  12.610 1.060 13.190 1.310 ;
        RECT  12.610 1.060 12.850 2.610 ;
        RECT  12.740 2.370 12.980 3.500 ;
        RECT  12.410 3.230 12.980 3.500 ;
        RECT  13.230 2.450 13.760 2.850 ;
        RECT  12.130 0.980 12.370 2.990 ;
        RECT  11.750 2.750 12.370 2.990 ;
        RECT  11.750 2.750 11.990 3.980 ;
        RECT  13.230 2.450 13.470 3.980 ;
        RECT  11.750 3.740 13.470 3.980 ;
        RECT  14.340 1.210 14.600 1.820 ;
        RECT  13.110 1.580 15.050 1.820 ;
        RECT  13.110 1.580 13.370 2.140 ;
        RECT  14.790 1.580 15.050 2.470 ;
        RECT  14.000 1.580 14.240 3.540 ;
        RECT  13.710 3.140 14.240 3.540 ;
        RECT  15.250 3.710 16.730 3.960 ;
        RECT  16.490 1.030 16.730 3.960 ;
        RECT  9.660 3.750 11.240 3.990 ;
        RECT  13.710 3.790 15.500 4.040 ;
        RECT  11.000 3.750 11.240 4.470 ;
        RECT  13.710 3.790 13.950 4.470 ;
        RECT  11.000 4.230 13.950 4.470 ;
        RECT  9.660 3.750 9.900 4.620 ;
        RECT  9.080 4.380 9.900 4.620 ;
        RECT  17.970 1.210 18.230 1.920 ;
        RECT  16.970 1.680 18.230 1.920 ;
        RECT  16.970 1.680 17.210 3.590 ;
        RECT  16.970 3.190 17.380 3.590 ;
    END
END slnht1

MACRO slnhq4
    CLASS CORE ;
    FOREIGN slnhq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.660 2.210 4.350 2.450 ;
        RECT  3.950 2.050 4.350 2.450 ;
        RECT  3.420 2.580 3.920 3.020 ;
        RECT  3.660 2.210 3.920 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.540 2.410 18.920 3.610 ;
        RECT  18.120 2.410 18.920 3.120 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.837  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.170 1.480 9.200 1.720 ;
        RECT  8.960 1.070 9.200 1.720 ;
        RECT  7.570 2.590 8.910 2.830 ;
        RECT  7.170 1.480 7.780 2.810 ;
        RECT  7.480 1.080 7.720 2.810 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        RECT  1.970 2.450 2.740 2.690 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.833  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.910 1.510 15.150 2.120 ;
        RECT  13.170 1.880 15.150 2.120 ;
        RECT  12.840 2.930 14.720 3.330 ;
        RECT  13.430 1.520 13.670 2.120 ;
        RECT  12.840 1.920 13.380 3.330 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.040 5.600 ;
        RECT  17.540 4.400 17.940 5.600 ;
        RECT  15.030 4.400 15.430 5.600 ;
        RECT  13.720 4.400 14.120 5.600 ;
        RECT  12.240 4.400 12.640 5.600 ;
        RECT  9.060 4.040 9.640 4.280 ;
        RECT  9.060 4.040 9.300 5.600 ;
        RECT  7.760 4.040 8.320 4.280 ;
        RECT  7.760 4.040 8.000 5.600 ;
        RECT  6.270 4.040 6.830 4.280 ;
        RECT  6.270 4.040 6.510 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.800 3.550 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.040 0.740 ;
        RECT  17.780 0.000 18.180 1.090 ;
        RECT  15.650 0.000 15.890 1.640 ;
        RECT  14.090 0.000 14.490 1.640 ;
        RECT  12.610 0.000 13.010 1.640 ;
        RECT  9.620 0.000 10.020 1.240 ;
        RECT  8.140 0.000 8.540 1.200 ;
        RECT  6.660 0.000 7.060 1.200 ;
        RECT  3.240 0.000 3.640 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.430 1.220 1.670 ;
        RECT  0.980 1.430 1.220 3.310 ;
        RECT  0.980 2.520 1.250 2.940 ;
        RECT  0.980 2.520 1.230 3.310 ;
        RECT  0.230 3.070 1.230 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.510 1.620 1.910 2.180 ;
        RECT  1.510 1.940 3.390 2.160 ;
        RECT  2.360 1.920 3.390 2.160 ;
        RECT  1.490 2.030 2.600 2.180 ;
        RECT  1.510 1.620 1.730 3.210 ;
        RECT  1.490 2.030 1.520 4.620 ;
        RECT  1.470 3.040 1.710 3.840 ;
        RECT  1.280 4.360 1.860 4.600 ;
        RECT  1.280 3.600 1.520 4.620 ;
        RECT  2.040 1.010 2.840 1.250 ;
        RECT  2.600 1.010 2.840 1.680 ;
        RECT  4.440 1.050 4.830 1.680 ;
        RECT  2.600 1.440 4.830 1.680 ;
        RECT  4.590 1.050 4.830 3.050 ;
        RECT  4.290 2.810 4.610 3.670 ;
        RECT  4.210 3.220 4.610 3.670 ;
        RECT  2.070 3.430 4.610 3.670 ;
        RECT  2.070 3.430 2.310 3.990 ;
        RECT  5.740 1.150 6.320 1.390 ;
        RECT  5.740 1.150 5.980 3.100 ;
        RECT  10.440 0.980 10.680 1.720 ;
        RECT  9.440 1.480 10.680 1.720 ;
        RECT  6.220 1.730 6.460 3.320 ;
        RECT  9.440 1.480 9.680 3.320 ;
        RECT  6.220 3.080 10.360 3.320 ;
        RECT  9.930 1.960 10.180 2.840 ;
        RECT  9.930 2.540 10.860 2.840 ;
        RECT  5.260 1.070 5.500 3.800 ;
        RECT  10.620 2.540 10.860 3.800 ;
        RECT  5.030 3.560 10.860 3.800 ;
        RECT  5.030 3.560 5.270 4.270 ;
        RECT  11.650 1.520 12.270 1.760 ;
        RECT  11.650 1.520 11.890 3.110 ;
        RECT  11.580 2.860 11.820 3.540 ;
        RECT  10.920 1.060 11.500 1.300 ;
        RECT  10.920 1.060 11.160 1.980 ;
        RECT  15.890 2.490 16.570 2.730 ;
        RECT  11.100 1.670 11.340 4.280 ;
        RECT  11.100 3.920 16.570 4.160 ;
        RECT  16.330 2.490 16.570 4.160 ;
        RECT  10.730 4.040 11.360 4.280 ;
        RECT  16.140 1.510 16.710 1.750 ;
        RECT  16.140 1.510 16.380 2.160 ;
        RECT  15.390 1.920 16.380 2.160 ;
        RECT  14.730 2.360 15.630 2.600 ;
        RECT  15.390 1.920 15.630 3.340 ;
        RECT  15.390 3.100 16.090 3.340 ;
        RECT  15.850 3.100 16.090 3.680 ;
        RECT  16.670 0.980 17.180 1.220 ;
        RECT  17.090 0.990 17.330 2.220 ;
        RECT  16.810 1.980 17.330 2.220 ;
        RECT  16.810 1.980 17.050 4.620 ;
        RECT  17.570 1.730 18.770 1.970 ;
        RECT  17.570 1.730 17.810 2.870 ;
        RECT  17.310 2.470 17.810 2.870 ;
        RECT  17.310 2.470 17.550 4.160 ;
        RECT  18.430 3.910 18.690 4.160 ;
        RECT  17.310 3.920 18.690 4.160 ;
        RECT  18.450 3.910 18.690 4.470 ;
    END
END slnhq4

MACRO slnhq2
    CLASS CORE ;
    FOREIGN slnhq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.660 2.210 4.350 2.450 ;
        RECT  3.950 2.050 4.350 2.450 ;
        RECT  3.420 2.580 3.920 3.020 ;
        RECT  3.660 2.210 3.920 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.900 16.120 3.610 ;
        RECT  15.290 2.900 16.120 3.140 ;
        RECT  15.290 2.430 15.530 3.140 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.980 1.480 7.720 1.720 ;
        RECT  7.480 1.070 7.720 1.720 ;
        RECT  6.980 2.590 7.680 2.830 ;
        RECT  6.980 1.480 7.220 2.830 ;
        RECT  6.780 2.020 7.220 2.460 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        RECT  1.970 2.450 2.740 2.690 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.260 1.920 12.190 2.160 ;
        RECT  11.950 1.510 12.190 2.160 ;
        RECT  11.460 3.010 12.150 3.250 ;
        RECT  11.460 1.920 11.700 3.250 ;
        RECT  11.260 1.920 11.700 2.460 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  14.790 4.400 15.190 5.600 ;
        RECT  12.350 4.400 12.750 5.600 ;
        RECT  10.830 4.400 11.230 5.600 ;
        RECT  7.720 4.040 8.280 4.280 ;
        RECT  7.720 4.040 7.960 5.600 ;
        RECT  6.200 4.040 6.760 4.280 ;
        RECT  6.200 4.040 6.440 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.800 3.550 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  14.820 0.000 15.220 1.090 ;
        RECT  12.690 0.000 12.930 1.640 ;
        RECT  11.130 0.000 11.530 1.640 ;
        RECT  8.140 0.000 8.540 1.200 ;
        RECT  6.660 0.000 7.060 1.200 ;
        RECT  3.240 0.000 3.640 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.430 1.220 1.670 ;
        RECT  0.980 1.430 1.220 3.310 ;
        RECT  0.980 2.520 1.250 2.940 ;
        RECT  0.930 2.930 1.230 3.310 ;
        RECT  0.230 3.070 1.230 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.490 1.620 1.910 2.170 ;
        RECT  1.490 1.930 3.390 2.170 ;
        RECT  2.990 1.930 3.390 2.330 ;
        RECT  1.490 1.620 1.730 3.190 ;
        RECT  1.470 3.040 1.710 3.840 ;
        RECT  1.280 4.360 1.860 4.600 ;
        RECT  1.280 3.600 1.520 4.620 ;
        RECT  2.040 1.010 2.850 1.250 ;
        RECT  2.610 1.010 2.850 1.680 ;
        RECT  4.440 1.050 4.830 1.680 ;
        RECT  2.610 1.440 4.830 1.680 ;
        RECT  4.200 3.200 4.830 3.670 ;
        RECT  4.590 1.050 4.830 3.670 ;
        RECT  2.070 3.430 4.830 3.670 ;
        RECT  2.070 3.430 2.310 3.990 ;
        RECT  5.740 1.150 6.320 1.390 ;
        RECT  5.740 1.150 6.000 3.100 ;
        RECT  5.740 2.780 6.010 3.100 ;
        RECT  8.960 0.980 9.200 1.720 ;
        RECT  7.960 1.480 9.200 1.720 ;
        RECT  7.960 2.740 9.020 2.980 ;
        RECT  6.250 1.740 6.490 3.320 ;
        RECT  7.960 1.480 8.200 3.320 ;
        RECT  6.250 3.080 8.200 3.320 ;
        RECT  8.460 1.960 8.700 2.500 ;
        RECT  8.460 2.260 9.500 2.500 ;
        RECT  9.260 2.260 9.500 3.460 ;
        RECT  8.770 3.220 9.500 3.460 ;
        RECT  8.770 3.220 9.010 3.800 ;
        RECT  5.260 3.560 9.010 3.800 ;
        RECT  5.260 1.070 5.500 4.190 ;
        RECT  4.950 3.950 5.500 4.190 ;
        RECT  10.240 1.520 10.790 1.760 ;
        RECT  10.240 1.520 10.480 3.540 ;
        RECT  13.180 1.510 13.750 1.750 ;
        RECT  13.180 1.510 13.420 2.160 ;
        RECT  12.430 1.920 13.420 2.160 ;
        RECT  12.040 2.480 12.670 2.720 ;
        RECT  12.430 1.920 12.670 3.680 ;
        RECT  13.170 3.100 13.410 3.680 ;
        RECT  12.430 3.440 13.410 3.680 ;
        RECT  9.620 0.980 9.980 1.380 ;
        RECT  12.930 2.410 13.330 2.860 ;
        RECT  12.930 2.620 13.890 2.860 ;
        RECT  9.740 0.980 9.980 4.160 ;
        RECT  9.390 3.840 9.980 4.080 ;
        RECT  13.650 2.620 13.890 4.160 ;
        RECT  9.740 3.920 13.890 4.160 ;
        RECT  13.710 0.980 14.370 1.220 ;
        RECT  14.130 0.980 14.370 4.620 ;
        RECT  14.610 1.730 15.810 1.970 ;
        RECT  14.610 1.730 14.850 4.160 ;
        RECT  15.750 3.910 16.010 4.160 ;
        RECT  14.610 3.920 16.010 4.160 ;
        RECT  15.770 3.910 16.010 4.470 ;
    END
END slnhq2

MACRO slnhq1
    CLASS CORE ;
    FOREIGN slnhq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.030 2.050 4.270 2.600 ;
        RECT  3.660 2.360 4.270 2.600 ;
        RECT  3.420 2.580 3.920 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.380 2.200 13.160 2.600 ;
        RECT  12.380 2.190 12.820 3.020 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.265  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.660 1.740 8.340 2.460 ;
        RECT  7.880 0.980 8.120 2.460 ;
        RECT  7.660 1.740 7.900 2.910 ;
        RECT  7.540 0.980 8.120 1.220 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        RECT  1.980 2.450 2.740 2.690 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.670  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.170 2.580 15.560 3.020 ;
        RECT  15.210 2.580 15.450 4.220 ;
        RECT  15.170 1.770 15.410 3.700 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.680 5.600 ;
        RECT  14.410 4.620 14.810 5.600 ;
        RECT  13.060 4.400 13.460 5.600 ;
        RECT  11.050 4.400 11.450 5.600 ;
        RECT  8.140 3.730 8.540 5.600 ;
        RECT  6.370 3.960 6.610 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.800 3.550 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.680 0.740 ;
        RECT  14.240 0.000 14.640 0.980 ;
        RECT  13.350 0.000 13.770 0.980 ;
        RECT  11.410 0.000 11.650 1.640 ;
        RECT  8.360 0.000 8.600 1.320 ;
        RECT  6.660 0.000 7.060 1.200 ;
        RECT  3.240 0.000 3.640 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.430 1.250 1.670 ;
        RECT  1.010 1.430 1.250 3.310 ;
        RECT  0.230 3.070 1.250 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.590 1.620 1.830 2.170 ;
        RECT  1.590 1.930 3.400 2.170 ;
        RECT  1.490 1.940 1.730 3.840 ;
        RECT  1.280 3.600 1.520 4.600 ;
        RECT  1.280 4.360 1.860 4.600 ;
        RECT  2.040 1.010 2.710 1.250 ;
        RECT  2.470 1.010 2.710 1.680 ;
        RECT  4.520 1.050 4.760 1.680 ;
        RECT  2.470 1.440 4.760 1.680 ;
        RECT  4.520 1.050 4.750 3.100 ;
        RECT  4.510 1.440 4.530 3.820 ;
        RECT  4.290 2.860 4.530 3.820 ;
        RECT  2.070 3.390 2.810 3.630 ;
        RECT  2.560 3.580 4.530 3.820 ;
        RECT  2.070 3.390 2.310 4.000 ;
        RECT  5.770 1.150 6.320 1.390 ;
        RECT  5.770 1.150 6.010 3.100 ;
        RECT  6.580 1.460 7.420 1.700 ;
        RECT  6.350 1.640 6.820 1.880 ;
        RECT  5.260 1.070 5.500 2.600 ;
        RECT  6.350 1.640 6.590 3.710 ;
        RECT  5.030 3.470 6.600 3.710 ;
        RECT  5.030 2.310 5.270 4.270 ;
        RECT  8.840 0.980 9.420 1.220 ;
        RECT  6.940 2.140 7.180 3.390 ;
        RECT  8.840 0.980 9.080 3.390 ;
        RECT  6.940 3.150 9.200 3.390 ;
        RECT  8.960 3.150 9.200 4.300 ;
        RECT  10.320 1.790 10.560 2.360 ;
        RECT  10.190 2.120 10.430 4.080 ;
        RECT  10.190 3.840 10.760 4.080 ;
        RECT  9.700 0.980 11.170 1.220 ;
        RECT  10.930 0.980 11.170 2.120 ;
        RECT  10.930 1.880 11.660 2.120 ;
        RECT  11.420 1.880 11.660 2.890 ;
        RECT  9.700 0.980 9.940 4.300 ;
        RECT  12.770 1.700 13.840 1.940 ;
        RECT  13.510 2.610 13.930 3.030 ;
        RECT  13.600 1.700 13.840 3.080 ;
        RECT  13.220 2.840 13.840 3.080 ;
        RECT  13.220 2.840 13.470 3.510 ;
        RECT  12.400 3.270 13.470 3.510 ;
        RECT  12.430 0.980 13.020 1.220 ;
        RECT  12.750 1.220 14.450 1.460 ;
        RECT  14.210 1.220 14.450 3.560 ;
        RECT  13.710 3.320 14.450 3.560 ;
        RECT  11.900 1.580 12.470 1.820 ;
        RECT  10.710 2.560 10.950 3.600 ;
        RECT  11.900 1.580 12.140 3.600 ;
        RECT  10.710 3.360 12.140 3.600 ;
        RECT  11.550 3.360 11.790 4.080 ;
        RECT  14.690 2.300 14.930 4.080 ;
        RECT  11.550 3.840 14.930 4.080 ;
    END
END slnhq1

MACRO slnhn4
    CLASS CORE ;
    FOREIGN slnhn4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.650 1.820 5.050 2.220 ;
        RECT  4.540 2.020 4.980 2.460 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.370 2.090 5.810 2.490 ;
        RECT  4.540 2.700 5.610 2.940 ;
        RECT  5.370 2.090 5.610 2.940 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.540 3.700 5.540 3.940 ;
        RECT  4.540 2.700 4.780 3.940 ;
        END
    END E
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.567  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.540 1.610 11.980 2.010 ;
        RECT  9.540 3.720 11.740 4.120 ;
        RECT  9.540 2.580 10.020 3.020 ;
        RECT  9.540 1.610 9.940 4.120 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.480 0.620 2.880 ;
        RECT  0.120 2.480 0.490 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.440 3.410 2.840 ;
        RECT  2.860 2.020 3.300 2.840 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.760  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.940 2.580 19.480 3.020 ;
        RECT  18.940 1.450 19.380 3.020 ;
        RECT  17.000 3.560 19.340 3.960 ;
        RECT  18.940 1.450 19.340 3.960 ;
        RECT  17.500 1.620 19.380 2.020 ;
        RECT  17.500 1.450 17.980 2.020 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.600 5.600 ;
        RECT  19.120 4.450 19.360 5.600 ;
        RECT  17.670 4.450 17.910 5.600 ;
        RECT  16.320 4.450 16.560 5.600 ;
        RECT  14.950 4.150 15.190 5.600 ;
        RECT  12.070 4.360 12.310 5.600 ;
        RECT  10.690 4.360 10.930 5.600 ;
        RECT  9.350 4.360 9.590 5.600 ;
        RECT  5.880 3.760 6.120 5.600 ;
        RECT  4.400 4.400 4.800 5.600 ;
        RECT  2.180 4.400 2.580 5.600 ;
        RECT  0.970 4.100 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.600 0.740 ;
        RECT  18.320 0.000 18.560 1.350 ;
        RECT  16.840 0.000 17.080 1.350 ;
        RECT  15.190 0.000 15.590 1.020 ;
        RECT  12.170 0.000 12.570 0.890 ;
        RECT  10.810 0.000 11.210 0.890 ;
        RECT  5.510 0.000 5.910 0.890 ;
        RECT  4.490 0.000 4.890 0.890 ;
        RECT  1.750 0.000 2.130 1.200 ;
        RECT  0.150 0.000 0.550 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.100 2.090 ;
        RECT  0.860 2.520 1.510 2.920 ;
        RECT  0.860 1.850 1.100 3.500 ;
        RECT  0.150 3.260 1.100 3.500 ;
        RECT  1.510 1.500 1.990 1.900 ;
        RECT  3.900 2.200 4.300 2.600 ;
        RECT  1.750 1.500 1.990 3.910 ;
        RECT  1.480 3.420 1.990 3.910 ;
        RECT  3.900 2.200 4.140 3.910 ;
        RECT  1.480 3.670 4.140 3.910 ;
        RECT  5.290 1.610 6.290 1.850 ;
        RECT  6.050 2.250 6.660 2.650 ;
        RECT  6.050 1.610 6.290 3.420 ;
        RECT  5.200 3.180 6.290 3.420 ;
        RECT  6.650 1.460 7.050 2.010 ;
        RECT  6.900 2.240 7.350 2.640 ;
        RECT  6.900 1.770 7.140 3.300 ;
        RECT  6.530 2.900 7.140 3.300 ;
        RECT  6.140 0.980 7.930 1.220 ;
        RECT  2.370 1.130 6.370 1.370 ;
        RECT  3.260 1.050 3.660 1.460 ;
        RECT  7.350 0.980 7.930 1.550 ;
        RECT  7.690 0.980 7.930 3.120 ;
        RECT  7.380 2.880 7.930 3.120 ;
        RECT  2.370 1.130 2.610 3.420 ;
        RECT  2.370 3.180 3.660 3.420 ;
        RECT  7.380 2.880 7.620 4.300 ;
        RECT  7.080 3.900 7.620 4.300 ;
        RECT  8.860 1.530 9.260 1.930 ;
        RECT  8.650 3.730 9.150 3.970 ;
        RECT  8.910 1.530 9.150 3.970 ;
        RECT  8.530 3.970 8.930 4.370 ;
        RECT  8.200 0.980 10.570 1.220 ;
        RECT  10.330 1.130 12.570 1.370 ;
        RECT  8.200 0.980 8.440 1.970 ;
        RECT  12.330 1.130 12.570 2.850 ;
        RECT  12.330 2.450 12.880 2.850 ;
        RECT  8.170 1.660 8.410 3.760 ;
        RECT  7.880 3.360 8.410 3.760 ;
        RECT  12.860 1.030 13.360 1.430 ;
        RECT  10.270 2.260 11.660 2.660 ;
        RECT  10.270 2.260 10.670 3.390 ;
        RECT  13.120 1.030 13.360 3.390 ;
        RECT  10.270 3.150 13.360 3.390 ;
        RECT  14.500 1.040 14.740 1.950 ;
        RECT  14.080 1.710 14.740 1.950 ;
        RECT  14.080 1.710 14.320 3.230 ;
        RECT  14.080 2.830 14.670 3.230 ;
        RECT  13.600 1.040 14.100 1.440 ;
        RECT  15.460 1.980 15.860 2.380 ;
        RECT  15.460 1.980 15.700 3.070 ;
        RECT  14.920 2.830 15.700 3.070 ;
        RECT  13.600 1.040 13.840 4.050 ;
        RECT  13.600 3.470 15.160 3.710 ;
        RECT  14.920 2.830 15.160 3.710 ;
        RECT  13.500 3.650 13.920 4.050 ;
        RECT  15.850 1.270 16.360 1.740 ;
        RECT  14.980 1.500 16.360 1.740 ;
        RECT  14.980 1.500 15.220 2.590 ;
        RECT  14.560 2.190 15.220 2.590 ;
        RECT  16.100 2.520 18.530 2.920 ;
        RECT  16.100 1.270 16.340 3.630 ;
        RECT  15.630 3.310 16.340 3.630 ;
    END
END slnhn4

MACRO slnhn2
    CLASS CORE ;
    FOREIGN slnhn2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.650 1.820 5.050 2.220 ;
        RECT  4.540 2.020 4.980 2.460 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.370 2.090 5.810 2.490 ;
        RECT  4.540 2.700 5.610 2.940 ;
        RECT  5.370 2.090 5.610 2.940 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.540 3.700 5.540 3.940 ;
        RECT  4.540 2.700 4.780 3.940 ;
        END
    END E
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.549  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.540 1.630 10.620 1.870 ;
        RECT  9.540 3.660 10.320 4.060 ;
        RECT  9.540 2.580 10.020 3.020 ;
        RECT  9.540 1.630 9.940 4.060 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.480 0.620 2.880 ;
        RECT  0.120 2.480 0.490 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.440 3.410 2.840 ;
        RECT  2.860 2.020 3.300 2.840 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.593  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.170 2.580 16.680 3.020 ;
        RECT  16.170 1.710 16.540 3.020 ;
        RECT  15.680 3.140 16.410 3.380 ;
        RECT  16.170 1.710 16.410 3.380 ;
        RECT  16.140 1.710 16.540 2.110 ;
        RECT  15.680 3.140 15.920 4.040 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  16.280 4.450 16.520 5.600 ;
        RECT  14.940 4.450 15.180 5.600 ;
        RECT  13.550 4.150 13.790 5.600 ;
        RECT  10.650 4.360 10.890 5.600 ;
        RECT  9.350 4.360 9.590 5.600 ;
        RECT  5.870 3.770 6.110 5.600 ;
        RECT  4.400 4.400 4.800 5.600 ;
        RECT  2.180 4.400 2.580 5.600 ;
        RECT  0.970 4.100 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  15.480 0.000 15.720 1.150 ;
        RECT  13.830 0.000 14.230 1.020 ;
        RECT  10.810 0.000 11.210 0.890 ;
        RECT  5.510 0.000 5.910 0.890 ;
        RECT  4.490 0.000 4.890 0.890 ;
        RECT  1.750 0.000 2.130 1.200 ;
        RECT  0.150 0.000 0.550 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.100 2.090 ;
        RECT  0.860 2.520 1.510 2.920 ;
        RECT  0.860 1.850 1.100 3.500 ;
        RECT  0.150 3.260 1.100 3.500 ;
        RECT  1.510 1.500 1.990 1.900 ;
        RECT  3.900 2.200 4.300 2.600 ;
        RECT  1.750 1.500 1.990 3.910 ;
        RECT  1.480 3.420 1.990 3.910 ;
        RECT  3.900 2.200 4.140 3.910 ;
        RECT  1.480 3.670 4.140 3.910 ;
        RECT  5.290 1.610 6.290 1.850 ;
        RECT  6.050 2.280 6.660 2.680 ;
        RECT  6.050 1.610 6.290 3.420 ;
        RECT  5.200 3.180 6.290 3.420 ;
        RECT  6.730 1.460 6.970 2.040 ;
        RECT  6.900 2.230 7.350 2.630 ;
        RECT  6.900 1.810 7.140 3.320 ;
        RECT  6.530 2.920 7.140 3.320 ;
        RECT  6.140 0.980 7.830 1.220 ;
        RECT  2.370 1.130 6.370 1.370 ;
        RECT  7.350 0.980 7.830 1.550 ;
        RECT  7.590 0.980 7.830 3.120 ;
        RECT  2.370 1.130 2.610 3.420 ;
        RECT  2.370 3.180 3.660 3.420 ;
        RECT  7.380 2.880 7.620 4.450 ;
        RECT  7.080 4.050 7.620 4.450 ;
        RECT  8.860 1.550 9.260 1.950 ;
        RECT  8.650 3.730 9.150 4.050 ;
        RECT  8.910 1.550 9.150 4.050 ;
        RECT  8.510 4.050 8.910 4.450 ;
        RECT  8.200 0.980 9.800 1.220 ;
        RECT  9.560 1.130 11.220 1.370 ;
        RECT  8.200 0.980 8.440 1.970 ;
        RECT  10.980 1.130 11.220 2.850 ;
        RECT  10.980 2.450 11.520 2.850 ;
        RECT  8.170 1.520 8.410 3.760 ;
        RECT  7.880 3.360 8.410 3.760 ;
        RECT  11.580 1.030 12.000 1.430 ;
        RECT  10.350 2.280 10.590 3.390 ;
        RECT  11.760 1.030 12.000 3.390 ;
        RECT  10.350 3.150 12.000 3.390 ;
        RECT  13.140 1.040 13.380 1.950 ;
        RECT  12.740 1.710 13.380 1.950 ;
        RECT  12.740 1.710 12.980 3.230 ;
        RECT  12.740 2.830 13.270 3.230 ;
        RECT  12.260 1.040 12.720 1.440 ;
        RECT  14.380 1.980 14.780 2.380 ;
        RECT  14.540 1.980 14.780 3.070 ;
        RECT  13.560 2.830 14.780 3.070 ;
        RECT  12.260 3.470 13.800 3.710 ;
        RECT  13.560 2.830 13.800 3.710 ;
        RECT  12.260 1.040 12.500 4.020 ;
        RECT  12.100 3.620 12.500 4.020 ;
        RECT  14.600 1.270 15.000 1.740 ;
        RECT  13.620 1.500 15.440 1.740 ;
        RECT  13.620 1.500 13.860 2.590 ;
        RECT  13.220 2.190 13.860 2.590 ;
        RECT  15.200 2.460 15.930 2.860 ;
        RECT  15.200 1.500 15.440 3.550 ;
        RECT  14.210 3.310 15.440 3.550 ;
    END
END slnhn2

MACRO slnhn1
    CLASS CORE ;
    FOREIGN slnhn1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.650 1.820 5.050 2.220 ;
        RECT  4.540 2.020 4.980 2.460 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.370 2.240 5.810 2.640 ;
        RECT  4.540 2.700 5.610 2.940 ;
        RECT  5.370 2.240 5.610 2.940 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.540 3.700 5.540 3.940 ;
        RECT  4.540 2.700 4.780 3.940 ;
        END
    END E
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.218  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.500 1.630 10.520 1.870 ;
        RECT  9.340 3.660 10.260 4.060 ;
        RECT  9.580 3.660 10.040 4.140 ;
        RECT  9.340 2.170 9.740 4.060 ;
        RECT  9.500 1.630 9.740 4.060 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.480 0.620 2.880 ;
        RECT  0.120 2.480 0.490 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.440 3.410 2.840 ;
        RECT  2.860 2.020 3.300 2.840 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.228  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.600 3.970 16.120 4.370 ;
        RECT  15.800 1.460 16.120 4.370 ;
        RECT  15.740 1.460 16.120 2.180 ;
        RECT  15.100 1.520 16.120 1.760 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  14.850 4.450 15.250 5.600 ;
        RECT  13.320 4.350 13.720 5.600 ;
        RECT  10.560 4.360 10.960 5.600 ;
        RECT  9.270 4.400 9.670 5.600 ;
        RECT  5.790 3.920 6.190 5.600 ;
        RECT  4.400 4.400 4.800 5.600 ;
        RECT  2.180 4.400 2.580 5.600 ;
        RECT  0.890 4.100 1.290 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  15.620 0.000 16.020 1.090 ;
        RECT  12.280 0.000 12.680 0.890 ;
        RECT  10.640 0.000 11.040 0.890 ;
        RECT  5.510 0.000 5.910 0.890 ;
        RECT  4.490 0.000 4.890 0.890 ;
        RECT  1.750 0.000 2.130 1.200 ;
        RECT  0.150 0.000 0.550 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.100 2.090 ;
        RECT  0.860 2.520 1.510 2.920 ;
        RECT  0.860 1.850 1.100 3.500 ;
        RECT  0.150 3.260 1.100 3.500 ;
        RECT  1.510 1.500 1.990 1.900 ;
        RECT  3.900 2.200 4.300 2.600 ;
        RECT  1.750 1.500 1.990 3.910 ;
        RECT  1.480 3.420 1.990 3.910 ;
        RECT  3.900 2.200 4.140 3.910 ;
        RECT  1.480 3.670 4.140 3.910 ;
        RECT  5.290 1.610 6.290 1.850 ;
        RECT  6.050 2.390 6.620 2.790 ;
        RECT  6.050 1.610 6.290 3.420 ;
        RECT  5.200 3.180 6.290 3.420 ;
        RECT  6.650 1.680 7.140 2.080 ;
        RECT  6.900 2.240 7.320 2.640 ;
        RECT  6.900 1.680 7.140 3.450 ;
        RECT  6.530 3.050 7.140 3.450 ;
        RECT  6.140 0.980 7.620 1.220 ;
        RECT  2.370 1.130 6.370 1.370 ;
        RECT  7.180 0.980 7.620 1.400 ;
        RECT  3.260 1.050 3.660 1.460 ;
        RECT  7.380 0.980 7.620 1.990 ;
        RECT  7.560 1.750 7.800 3.120 ;
        RECT  2.370 1.130 2.610 3.420 ;
        RECT  2.370 3.180 3.660 3.420 ;
        RECT  7.380 2.880 7.620 4.300 ;
        RECT  7.070 3.900 7.620 4.300 ;
        RECT  8.700 1.550 9.100 2.360 ;
        RECT  8.630 2.120 8.870 4.370 ;
        RECT  8.520 3.970 8.920 4.370 ;
        RECT  8.040 0.980 10.400 1.220 ;
        RECT  10.160 1.130 11.100 1.370 ;
        RECT  10.860 1.130 11.100 2.850 ;
        RECT  10.660 2.450 11.100 2.850 ;
        RECT  8.040 0.980 8.280 3.760 ;
        RECT  7.870 3.360 8.280 3.760 ;
        RECT  11.340 1.220 11.810 1.620 ;
        RECT  9.980 2.280 10.380 2.680 ;
        RECT  10.140 2.280 10.380 3.390 ;
        RECT  10.140 3.150 11.580 3.390 ;
        RECT  11.340 1.220 11.580 3.510 ;
        RECT  11.150 3.110 11.580 3.510 ;
        RECT  12.870 1.230 13.290 1.630 ;
        RECT  12.870 1.230 13.110 2.110 ;
        RECT  12.720 1.870 12.960 3.350 ;
        RECT  12.720 2.950 13.120 3.350 ;
        RECT  12.150 1.230 12.550 1.630 ;
        RECT  12.150 1.230 12.400 2.120 ;
        RECT  11.820 1.880 12.400 2.120 ;
        RECT  14.030 2.420 14.430 2.820 ;
        RECT  14.030 2.420 14.270 3.530 ;
        RECT  13.560 3.290 14.270 3.530 ;
        RECT  11.820 1.880 12.060 3.990 ;
        RECT  13.560 3.290 13.800 3.830 ;
        RECT  11.820 3.590 13.800 3.830 ;
        RECT  11.820 3.590 12.350 3.990 ;
        RECT  14.250 1.040 14.650 2.180 ;
        RECT  13.350 1.940 14.910 2.180 ;
        RECT  13.350 1.940 13.750 2.390 ;
        RECT  14.670 2.570 15.560 2.940 ;
        RECT  14.670 1.940 14.910 4.190 ;
        RECT  14.050 3.790 14.910 4.190 ;
    END
END slnhn1

MACRO slnhb4
    CLASS CORE ;
    FOREIGN slnhb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.660 2.210 4.350 2.460 ;
        RECT  3.950 2.040 4.350 2.460 ;
        RECT  3.420 2.580 3.920 3.020 ;
        RECT  3.660 2.210 3.920 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  21.280 2.020 21.720 2.460 ;
        RECT  21.020 2.310 21.540 2.550 ;
        RECT  21.020 2.310 21.420 2.710 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.724  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.440 1.480 12.160 1.720 ;
        RECT  11.920 1.070 12.160 1.720 ;
        RECT  10.530 2.590 11.940 2.830 ;
        RECT  10.130 2.570 11.140 2.810 ;
        RECT  10.700 1.480 11.140 2.830 ;
        RECT  10.440 1.080 10.680 1.720 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.146  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.710 1.150 9.280 1.390 ;
        RECT  6.880 2.590 8.980 2.830 ;
        RECT  7.170 1.480 8.960 1.720 ;
        RECT  8.710 1.150 8.960 1.720 ;
        RECT  7.170 1.480 7.780 2.830 ;
        RECT  7.480 1.080 7.720 2.830 ;
        RECT  6.880 2.480 7.570 2.900 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        RECT  1.980 2.450 2.740 2.690 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.806  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 1.920 18.070 2.160 ;
        RECT  17.830 1.510 18.070 2.160 ;
        RECT  15.740 3.010 17.690 3.250 ;
        RECT  16.350 1.520 16.590 2.160 ;
        RECT  15.950 1.920 16.350 3.330 ;
        RECT  15.740 1.920 16.350 3.250 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 21.840 5.600 ;
        RECT  20.380 3.450 20.950 3.690 ;
        RECT  20.380 3.450 20.620 5.600 ;
        RECT  18.000 4.400 18.400 5.600 ;
        RECT  16.340 4.400 16.740 5.600 ;
        RECT  15.040 4.400 15.440 5.600 ;
        RECT  12.030 4.040 12.630 4.280 ;
        RECT  12.030 4.040 12.270 5.600 ;
        RECT  10.260 4.040 10.930 4.280 ;
        RECT  10.260 4.040 10.500 5.600 ;
        RECT  9.060 4.040 9.670 4.280 ;
        RECT  9.060 4.040 9.300 5.600 ;
        RECT  7.760 4.040 8.360 4.280 ;
        RECT  7.760 4.040 8.000 5.600 ;
        RECT  6.250 4.040 6.870 4.280 ;
        RECT  6.250 4.040 6.490 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.800 3.550 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 21.840 0.740 ;
        RECT  20.540 0.000 20.990 1.030 ;
        RECT  18.570 0.000 18.810 1.640 ;
        RECT  17.090 0.000 17.330 1.640 ;
        RECT  15.610 0.000 15.850 1.640 ;
        RECT  12.660 0.000 12.900 1.240 ;
        RECT  11.100 0.000 11.500 1.240 ;
        RECT  9.620 0.000 10.020 1.200 ;
        RECT  8.220 0.000 8.460 1.240 ;
        RECT  6.660 0.000 7.060 1.200 ;
        RECT  3.240 0.000 3.640 1.200 ;
        RECT  0.730 0.000 1.150 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.140 1.430 1.260 1.670 ;
        RECT  1.020 1.430 1.260 3.310 ;
        RECT  0.230 3.070 1.260 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.500 1.620 1.920 2.170 ;
        RECT  1.500 1.930 3.400 2.170 ;
        RECT  1.500 1.620 1.740 3.840 ;
        RECT  1.280 4.360 1.860 4.600 ;
        RECT  1.280 3.600 1.520 4.620 ;
        RECT  2.040 1.010 2.780 1.250 ;
        RECT  2.540 1.010 2.780 1.680 ;
        RECT  4.440 1.050 4.840 1.680 ;
        RECT  2.540 1.440 4.840 1.680 ;
        RECT  4.180 3.160 4.840 3.820 ;
        RECT  2.070 3.420 3.630 3.660 ;
        RECT  4.600 1.050 4.840 3.820 ;
        RECT  3.290 3.580 4.840 3.820 ;
        RECT  2.070 3.420 2.310 4.000 ;
        RECT  5.740 1.150 6.320 1.390 ;
        RECT  5.740 1.150 5.980 2.180 ;
        RECT  5.620 1.880 5.860 3.100 ;
        RECT  13.160 0.980 13.720 1.220 ;
        RECT  13.160 0.980 13.400 1.720 ;
        RECT  12.400 1.480 13.400 1.720 ;
        RECT  9.160 1.900 9.740 2.140 ;
        RECT  12.400 1.480 12.640 3.320 ;
        RECT  9.500 1.900 9.740 3.320 ;
        RECT  12.400 2.740 12.650 3.320 ;
        RECT  9.500 3.080 13.340 3.320 ;
        RECT  5.260 1.070 5.500 1.640 ;
        RECT  12.900 1.960 13.150 2.650 ;
        RECT  12.900 2.410 13.820 2.650 ;
        RECT  5.080 1.400 5.320 3.800 ;
        RECT  13.580 2.410 13.820 3.800 ;
        RECT  5.080 3.560 13.820 3.800 ;
        RECT  5.370 3.560 5.610 4.430 ;
        RECT  4.940 4.190 5.610 4.430 ;
        RECT  14.620 1.690 14.860 3.540 ;
        RECT  14.460 3.130 14.880 3.540 ;
        RECT  14.060 0.980 15.360 1.220 ;
        RECT  18.830 2.470 19.540 2.710 ;
        RECT  15.120 0.980 15.360 4.160 ;
        RECT  14.060 3.920 19.540 4.160 ;
        RECT  19.300 2.470 19.540 4.160 ;
        RECT  13.690 4.040 14.300 4.280 ;
        RECT  19.060 1.510 19.640 1.750 ;
        RECT  19.060 1.510 19.300 2.160 ;
        RECT  18.350 1.920 19.300 2.160 ;
        RECT  17.670 2.480 18.590 2.720 ;
        RECT  18.350 1.920 18.590 3.340 ;
        RECT  18.350 3.100 19.060 3.340 ;
        RECT  18.820 3.100 19.060 3.680 ;
        RECT  19.590 0.980 20.250 1.220 ;
        RECT  20.010 0.980 20.250 2.220 ;
        RECT  19.780 1.980 20.020 3.660 ;
        RECT  20.530 1.510 21.690 1.750 ;
        RECT  20.530 1.510 20.770 2.700 ;
        RECT  20.260 2.460 20.770 2.700 ;
        RECT  20.260 2.460 20.500 3.210 ;
        RECT  20.260 2.970 21.610 3.210 ;
        RECT  21.370 2.970 21.610 3.550 ;
    END
END slnhb4

MACRO slnhb2
    CLASS CORE ;
    FOREIGN slnhb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.660 2.330 4.270 2.570 ;
        RECT  4.030 1.990 4.270 2.570 ;
        RECT  3.420 2.580 3.920 3.020 ;
        RECT  3.660 2.330 3.920 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.860 2.580 17.240 3.020 ;
        RECT  16.480 2.430 16.880 2.830 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.727  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 1.440 9.200 1.720 ;
        RECT  8.960 1.070 9.200 1.720 ;
        RECT  8.830 2.250 9.070 2.840 ;
        RECT  8.460 1.440 8.900 1.900 ;
        RECT  8.460 2.250 9.070 2.500 ;
        RECT  8.460 1.440 8.810 2.500 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.722  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.230 1.150 7.800 1.390 ;
        RECT  6.930 3.080 7.480 3.320 ;
        RECT  6.980 1.480 7.480 1.720 ;
        RECT  7.230 1.150 7.480 1.720 ;
        RECT  6.780 2.020 7.220 2.460 ;
        RECT  6.980 1.480 7.220 2.460 ;
        RECT  6.930 2.020 7.170 3.320 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        RECT  1.980 2.450 2.740 2.690 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.404  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.380 3.260 13.720 3.500 ;
        RECT  12.790 1.920 13.530 2.160 ;
        RECT  13.290 1.510 13.530 2.160 ;
        RECT  12.380 3.140 13.030 3.580 ;
        RECT  12.790 1.920 13.030 3.580 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.360 5.600 ;
        RECT  16.160 4.330 16.560 5.600 ;
        RECT  13.880 4.400 14.280 5.600 ;
        RECT  12.300 4.400 12.700 5.600 ;
        RECT  9.260 4.040 9.870 4.280 ;
        RECT  9.260 4.040 9.500 5.600 ;
        RECT  7.590 4.040 8.160 4.280 ;
        RECT  7.590 4.040 7.840 5.600 ;
        RECT  6.230 4.040 6.860 4.280 ;
        RECT  6.230 4.040 6.470 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.800 3.550 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.360 0.740 ;
        RECT  16.160 0.000 16.560 1.090 ;
        RECT  14.030 0.000 14.270 1.640 ;
        RECT  12.470 0.000 12.870 1.640 ;
        RECT  9.700 0.000 9.940 1.240 ;
        RECT  8.140 0.000 8.540 1.200 ;
        RECT  6.740 0.000 6.980 1.200 ;
        RECT  3.240 0.000 3.640 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.430 1.260 1.670 ;
        RECT  1.020 1.430 1.260 3.310 ;
        RECT  0.230 3.070 1.260 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.500 1.620 1.920 2.170 ;
        RECT  1.500 1.930 3.400 2.170 ;
        RECT  1.500 1.620 1.740 3.840 ;
        RECT  1.280 4.360 1.860 4.600 ;
        RECT  1.280 3.600 1.520 4.620 ;
        RECT  2.040 1.010 2.810 1.250 ;
        RECT  2.570 1.010 2.810 1.680 ;
        RECT  4.520 1.050 4.760 1.680 ;
        RECT  2.570 1.440 4.760 1.680 ;
        RECT  4.510 1.440 4.750 3.820 ;
        RECT  4.210 3.160 4.750 3.820 ;
        RECT  2.070 3.430 3.750 3.670 ;
        RECT  3.340 3.580 4.750 3.820 ;
        RECT  2.070 3.430 2.310 4.000 ;
        RECT  5.740 1.150 6.320 1.390 ;
        RECT  5.740 1.150 5.980 2.340 ;
        RECT  5.620 1.920 5.860 3.100 ;
        RECT  5.260 1.070 5.500 1.680 ;
        RECT  9.920 1.960 10.160 3.800 ;
        RECT  5.030 3.560 10.160 3.800 ;
        RECT  5.030 1.440 5.270 4.270 ;
        RECT  9.440 1.480 10.680 1.720 ;
        RECT  7.650 1.910 8.170 2.310 ;
        RECT  7.930 1.910 8.170 3.320 ;
        RECT  9.440 1.480 9.680 3.320 ;
        RECT  7.930 3.080 9.680 3.320 ;
        RECT  10.440 0.970 10.680 3.480 ;
        RECT  10.560 3.220 10.800 4.280 ;
        RECT  10.190 4.040 10.800 4.280 ;
        RECT  11.710 1.780 12.280 2.020 ;
        RECT  12.030 1.780 12.280 2.630 ;
        RECT  11.790 2.370 12.030 3.540 ;
        RECT  11.730 3.130 12.130 3.540 ;
        RECT  14.520 1.510 15.090 1.750 ;
        RECT  14.520 1.510 14.770 2.160 ;
        RECT  14.120 1.920 14.770 2.160 ;
        RECT  13.270 2.480 14.360 2.720 ;
        RECT  14.120 1.920 14.360 3.260 ;
        RECT  14.120 3.020 15.020 3.260 ;
        RECT  10.930 0.990 11.480 1.230 ;
        RECT  10.930 0.990 11.170 2.700 ;
        RECT  11.520 3.920 14.830 4.160 ;
        RECT  11.040 2.400 11.280 4.600 ;
        RECT  14.590 3.920 14.830 4.620 ;
        RECT  11.520 3.920 11.760 4.600 ;
        RECT  11.040 4.360 11.760 4.600 ;
        RECT  14.590 4.380 15.380 4.620 ;
        RECT  15.050 0.980 15.710 1.220 ;
        RECT  15.470 0.980 15.710 2.320 ;
        RECT  15.260 2.070 15.500 4.080 ;
        RECT  15.260 3.840 15.820 4.080 ;
        RECT  15.950 1.730 17.150 1.970 ;
        RECT  15.800 2.550 16.200 2.950 ;
        RECT  15.950 1.730 16.200 3.550 ;
        RECT  15.940 2.550 16.200 3.550 ;
        RECT  15.940 3.310 17.130 3.550 ;
    END
END slnhb2

MACRO slnhb1
    CLASS CORE ;
    FOREIGN slnhb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.660 2.210 4.360 2.450 ;
        RECT  3.420 2.580 3.920 3.020 ;
        RECT  3.660 2.210 3.920 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.940 2.300 13.420 3.020 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.110 2.020 8.900 2.460 ;
        RECT  8.180 1.510 8.440 2.460 ;
        RECT  8.180 1.090 8.420 2.460 ;
        RECT  8.110 1.770 8.350 2.890 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.261  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.600 1.440 7.720 1.680 ;
        RECT  7.480 1.090 7.720 1.680 ;
        RECT  6.500 3.080 7.290 3.320 ;
        RECT  6.220 2.020 6.840 2.460 ;
        RECT  6.600 1.440 6.840 2.460 ;
        RECT  6.500 2.020 6.740 3.320 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        RECT  1.980 2.450 2.740 2.690 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.715  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 1.460 16.120 1.900 ;
        RECT  15.770 1.460 16.010 4.530 ;
        RECT  15.740 1.460 16.010 1.920 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  14.960 4.620 15.360 5.600 ;
        RECT  13.610 4.400 14.010 5.600 ;
        RECT  11.590 4.400 11.990 5.600 ;
        RECT  8.410 3.980 9.070 4.220 ;
        RECT  8.410 3.980 8.650 5.600 ;
        RECT  6.130 4.040 6.760 4.280 ;
        RECT  6.130 4.040 6.370 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.800 3.550 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  14.820 0.000 15.250 0.980 ;
        RECT  13.950 0.000 14.370 0.980 ;
        RECT  12.010 0.000 12.250 1.640 ;
        RECT  8.920 0.000 9.160 1.320 ;
        RECT  6.660 0.000 7.060 1.200 ;
        RECT  3.240 0.000 3.640 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.430 1.260 1.670 ;
        RECT  0.990 1.430 1.260 2.940 ;
        RECT  0.940 2.930 1.230 3.310 ;
        RECT  0.230 3.070 1.230 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.500 1.620 1.920 2.170 ;
        RECT  1.500 1.930 3.400 2.170 ;
        RECT  1.480 3.170 1.740 3.840 ;
        RECT  1.500 1.620 1.740 3.840 ;
        RECT  1.280 4.360 1.860 4.600 ;
        RECT  1.280 3.600 1.520 4.620 ;
        RECT  2.040 1.010 2.760 1.250 ;
        RECT  2.520 1.010 2.760 1.680 ;
        RECT  4.400 1.050 4.870 1.680 ;
        RECT  2.520 1.440 4.870 1.680 ;
        RECT  4.630 1.050 4.870 3.320 ;
        RECT  4.210 2.980 4.790 3.820 ;
        RECT  2.070 3.430 3.330 3.670 ;
        RECT  2.980 3.580 4.790 3.820 ;
        RECT  2.070 3.430 2.310 4.000 ;
        RECT  5.740 1.150 6.320 1.390 ;
        RECT  5.740 1.150 5.980 2.130 ;
        RECT  5.620 1.870 5.860 3.100 ;
        RECT  5.260 1.070 5.500 1.630 ;
        RECT  5.120 1.390 5.360 3.800 ;
        RECT  5.030 3.560 7.340 3.800 ;
        RECT  7.100 3.560 7.340 4.500 ;
        RECT  5.030 3.560 5.270 4.270 ;
        RECT  7.100 4.260 7.860 4.500 ;
        RECT  9.410 0.980 9.980 1.220 ;
        RECT  7.630 1.960 7.870 3.370 ;
        RECT  9.410 0.980 9.650 3.370 ;
        RECT  7.630 3.130 9.740 3.370 ;
        RECT  9.500 3.130 9.740 4.300 ;
        RECT  10.790 1.790 11.290 2.320 ;
        RECT  10.790 1.790 11.030 3.380 ;
        RECT  10.730 3.060 10.970 4.080 ;
        RECT  10.730 3.840 11.300 4.080 ;
        RECT  10.240 0.980 11.770 1.220 ;
        RECT  11.530 0.980 11.770 2.120 ;
        RECT  11.530 1.880 12.200 2.120 ;
        RECT  11.960 1.880 12.200 2.970 ;
        RECT  10.240 0.980 10.480 4.300 ;
        RECT  13.370 1.700 14.420 1.940 ;
        RECT  14.170 1.700 14.420 3.080 ;
        RECT  14.170 2.440 14.570 3.080 ;
        RECT  13.740 2.840 14.570 3.080 ;
        RECT  13.740 2.840 13.980 3.600 ;
        RECT  12.960 3.360 13.980 3.600 ;
        RECT  13.030 0.980 13.670 1.220 ;
        RECT  13.420 1.220 15.050 1.460 ;
        RECT  14.810 1.220 15.050 3.560 ;
        RECT  14.260 3.320 15.050 3.560 ;
        RECT  12.750 1.500 12.990 2.060 ;
        RECT  12.440 1.810 12.990 2.060 ;
        RECT  11.270 2.560 11.510 3.600 ;
        RECT  12.440 1.810 12.680 3.600 ;
        RECT  11.270 3.360 12.680 3.600 ;
        RECT  12.010 3.360 12.250 4.080 ;
        RECT  15.290 2.290 15.530 4.080 ;
        RECT  12.010 3.840 15.530 4.080 ;
    END
END slnhb1

MACRO slclq4
    CLASS CORE ;
    FOREIGN slclq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.090 2.020 10.540 2.510 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.190 2.280 5.370 2.520 ;
        RECT  5.130 1.160 5.370 2.520 ;
        RECT  4.410 1.160 5.370 1.400 ;
        RECT  3.100 0.980 4.650 1.220 ;
        RECT  4.190 2.280 4.430 3.170 ;
        RECT  3.980 2.580 4.430 3.170 ;
        RECT  3.690 2.930 4.090 3.490 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.404  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 2.530 6.420 3.020 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.770  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.160 3.050 14.480 3.290 ;
        RECT  14.240 1.100 14.480 3.290 ;
        RECT  13.160 2.490 13.400 3.290 ;
        RECT  12.240 2.490 13.400 2.730 ;
        RECT  12.560 1.100 13.080 1.500 ;
        RECT  12.240 1.460 12.820 1.900 ;
        RECT  12.240 1.460 12.480 2.730 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.720 2.700 ;
        RECT  0.120 2.300 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.580 3.330 3.320 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.759  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.170 3.880 21.550 4.120 ;
        RECT  21.310 1.090 21.550 4.120 ;
        RECT  19.660 1.020 20.150 1.930 ;
        RECT  19.660 1.020 19.900 4.120 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 21.840 5.600 ;
        RECT  21.210 4.620 21.610 5.600 ;
        RECT  19.900 4.620 20.300 5.600 ;
        RECT  18.590 4.620 18.990 5.600 ;
        RECT  17.240 4.200 17.480 5.600 ;
        RECT  15.290 4.780 15.800 5.600 ;
        RECT  14.570 4.200 14.810 5.600 ;
        RECT  13.460 4.040 13.700 5.600 ;
        RECT  13.140 4.040 13.700 4.280 ;
        RECT  12.120 3.450 12.360 5.600 ;
        RECT  11.800 3.450 12.360 3.690 ;
        RECT  9.870 3.880 10.110 5.600 ;
        RECT  6.530 4.710 6.930 5.600 ;
        RECT  4.440 4.620 4.840 5.600 ;
        RECT  2.080 4.450 2.320 5.600 ;
        RECT  0.730 4.580 1.130 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 21.840 0.740 ;
        RECT  20.570 0.000 20.810 1.240 ;
        RECT  19.090 0.000 19.330 1.150 ;
        RECT  17.650 0.000 17.890 1.320 ;
        RECT  15.620 0.000 16.140 0.820 ;
        RECT  13.500 0.000 13.740 1.250 ;
        RECT  12.020 0.000 12.260 1.210 ;
        RECT  10.490 1.060 11.040 1.300 ;
        RECT  10.800 0.000 11.040 1.300 ;
        RECT  6.340 0.000 6.740 0.890 ;
        RECT  5.250 0.000 5.650 0.890 ;
        RECT  0.690 0.000 0.930 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.200 1.820 ;
        RECT  0.960 2.410 1.490 2.810 ;
        RECT  0.960 1.580 1.200 3.500 ;
        RECT  0.150 3.260 1.200 3.500 ;
        RECT  0.150 3.260 0.560 3.660 ;
        RECT  1.510 1.510 2.020 1.930 ;
        RECT  1.760 1.510 2.020 4.160 ;
        RECT  1.780 0.980 2.020 4.160 ;
        RECT  1.470 3.760 2.020 4.160 ;
        RECT  2.260 0.980 2.860 1.220 ;
        RECT  2.620 0.980 2.860 1.700 ;
        RECT  2.620 1.460 4.160 1.700 ;
        RECT  3.920 1.640 4.890 1.880 ;
        RECT  4.480 1.640 4.890 2.040 ;
        RECT  5.750 1.850 6.530 2.090 ;
        RECT  6.290 2.040 7.020 2.280 ;
        RECT  6.780 2.040 7.020 3.540 ;
        RECT  5.880 3.300 7.020 3.540 ;
        RECT  7.260 0.980 8.020 1.220 ;
        RECT  7.110 1.400 7.510 1.800 ;
        RECT  7.260 2.600 7.780 3.000 ;
        RECT  7.260 0.980 7.510 3.620 ;
        RECT  7.810 1.470 8.390 1.870 ;
        RECT  2.330 1.940 3.680 2.180 ;
        RECT  8.150 1.470 8.390 3.630 ;
        RECT  7.880 3.220 8.390 3.630 ;
        RECT  2.330 1.940 2.570 4.020 ;
        RECT  2.330 3.780 5.580 4.020 ;
        RECT  7.880 3.220 8.120 4.100 ;
        RECT  5.180 3.860 8.120 4.100 ;
        RECT  5.180 3.780 5.580 4.450 ;
        RECT  9.110 1.470 9.690 1.710 ;
        RECT  9.110 1.470 9.350 3.630 ;
        RECT  9.110 3.230 10.930 3.630 ;
        RECT  8.630 0.980 10.190 1.220 ;
        RECT  9.950 0.980 10.190 1.780 ;
        RECT  9.950 1.540 11.020 1.780 ;
        RECT  10.780 1.540 11.020 2.470 ;
        RECT  10.780 2.070 11.440 2.470 ;
        RECT  8.630 0.980 8.870 4.310 ;
        RECT  8.450 3.900 8.870 4.310 ;
        RECT  11.280 0.980 11.520 1.710 ;
        RECT  11.280 1.460 11.920 1.710 ;
        RECT  15.430 1.330 15.670 2.210 ;
        RECT  15.160 1.970 15.670 2.210 ;
        RECT  9.590 2.150 9.830 2.990 ;
        RECT  11.680 1.460 11.920 3.210 ;
        RECT  9.590 2.750 11.920 2.990 ;
        RECT  11.220 2.970 12.880 3.210 ;
        RECT  12.640 2.970 12.880 3.800 ;
        RECT  15.160 1.970 15.400 3.800 ;
        RECT  12.640 3.560 15.400 3.800 ;
        RECT  11.220 2.750 11.460 4.360 ;
        RECT  16.650 1.410 17.230 1.650 ;
        RECT  16.650 1.410 16.890 3.210 ;
        RECT  16.170 1.330 16.410 2.530 ;
        RECT  15.900 2.290 16.410 2.530 ;
        RECT  15.900 2.290 16.150 3.690 ;
        RECT  18.000 2.070 18.240 3.690 ;
        RECT  15.900 3.450 18.240 3.690 ;
        RECT  18.310 1.330 18.730 1.800 ;
        RECT  17.470 1.560 18.730 1.800 ;
        RECT  17.470 1.560 17.710 2.180 ;
        RECT  17.130 1.940 17.710 2.180 ;
        RECT  18.490 2.120 19.360 2.520 ;
        RECT  18.490 1.330 18.730 4.170 ;
        RECT  17.900 3.930 18.730 4.170 ;
    END
END slclq4

MACRO slclq2
    CLASS CORE ;
    FOREIGN slclq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.070 2.020 10.540 2.510 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.190 2.280 5.370 2.520 ;
        RECT  5.130 1.160 5.370 2.520 ;
        RECT  4.410 1.160 5.370 1.400 ;
        RECT  3.100 0.980 4.650 1.220 ;
        RECT  4.190 2.280 4.430 3.170 ;
        RECT  3.980 2.580 4.430 3.170 ;
        RECT  3.690 2.930 4.090 3.490 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.404  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 2.530 6.420 3.020 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.334  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.760 2.020 13.390 2.460 ;
        RECT  12.410 2.490 13.000 2.730 ;
        RECT  12.760 1.100 13.000 2.730 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.320 2.300 0.720 2.700 ;
        RECT  0.120 2.460 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.580 3.330 3.320 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.907  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.540 1.460 19.250 1.930 ;
        RECT  19.010 1.020 19.250 1.930 ;
        RECT  18.200 3.140 18.790 3.380 ;
        RECT  18.540 1.460 18.790 3.380 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.600 5.600 ;
        RECT  18.930 4.620 19.330 5.600 ;
        RECT  17.630 4.620 18.030 5.600 ;
        RECT  16.190 4.000 16.430 5.600 ;
        RECT  14.050 4.780 14.580 5.600 ;
        RECT  13.330 4.310 13.570 5.600 ;
        RECT  12.170 3.450 12.410 5.600 ;
        RECT  11.810 3.450 12.410 3.690 ;
        RECT  9.870 3.880 10.110 5.600 ;
        RECT  6.530 4.710 6.930 5.600 ;
        RECT  4.440 4.620 4.840 5.600 ;
        RECT  2.080 4.450 2.320 5.600 ;
        RECT  0.730 4.580 1.130 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.600 0.740 ;
        RECT  18.190 0.000 18.590 0.980 ;
        RECT  16.520 0.000 16.760 1.320 ;
        RECT  14.480 0.000 15.000 0.820 ;
        RECT  13.500 0.000 13.740 1.250 ;
        RECT  12.020 0.000 12.260 1.230 ;
        RECT  10.490 1.060 11.040 1.300 ;
        RECT  10.800 0.000 11.040 1.300 ;
        RECT  6.340 0.000 6.740 0.890 ;
        RECT  5.250 0.000 5.650 0.890 ;
        RECT  0.690 0.000 0.930 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.200 1.820 ;
        RECT  0.960 2.410 1.490 2.810 ;
        RECT  0.960 1.580 1.200 3.500 ;
        RECT  0.150 3.260 1.200 3.500 ;
        RECT  0.150 3.260 0.560 3.660 ;
        RECT  1.510 1.510 2.020 1.930 ;
        RECT  1.750 1.510 2.020 4.160 ;
        RECT  1.780 0.980 2.020 4.160 ;
        RECT  1.470 3.760 2.020 4.160 ;
        RECT  2.260 0.980 2.860 1.220 ;
        RECT  2.620 0.980 2.860 1.700 ;
        RECT  2.620 1.460 4.160 1.700 ;
        RECT  3.920 1.640 4.890 1.880 ;
        RECT  4.480 1.640 4.890 2.040 ;
        RECT  5.750 1.850 6.530 2.090 ;
        RECT  6.290 2.040 7.020 2.280 ;
        RECT  6.780 2.040 7.020 3.540 ;
        RECT  5.880 3.300 7.020 3.540 ;
        RECT  7.260 0.980 8.020 1.220 ;
        RECT  7.110 1.400 7.510 1.800 ;
        RECT  7.260 2.580 7.790 2.990 ;
        RECT  7.260 0.980 7.510 3.620 ;
        RECT  7.810 1.470 8.380 1.870 ;
        RECT  2.330 1.940 3.680 2.180 ;
        RECT  8.140 1.470 8.380 3.630 ;
        RECT  7.880 3.220 8.380 3.630 ;
        RECT  2.330 1.940 2.570 4.020 ;
        RECT  2.330 3.780 5.580 4.020 ;
        RECT  7.880 3.220 8.120 4.100 ;
        RECT  5.180 3.860 8.120 4.100 ;
        RECT  5.180 3.780 5.580 4.450 ;
        RECT  9.110 1.470 9.690 1.710 ;
        RECT  9.110 1.470 9.350 3.630 ;
        RECT  9.110 3.230 10.930 3.630 ;
        RECT  8.630 0.980 10.190 1.220 ;
        RECT  9.950 0.980 10.190 1.780 ;
        RECT  9.950 1.540 11.030 1.780 ;
        RECT  10.790 1.540 11.030 2.430 ;
        RECT  10.790 2.190 11.450 2.430 ;
        RECT  8.630 0.980 8.870 4.310 ;
        RECT  8.450 3.900 8.870 4.310 ;
        RECT  11.280 0.990 11.520 1.950 ;
        RECT  11.280 1.710 11.930 1.950 ;
        RECT  14.300 1.330 14.540 2.210 ;
        RECT  14.030 1.970 14.540 2.210 ;
        RECT  9.590 2.150 9.830 2.990 ;
        RECT  11.690 1.710 11.930 3.210 ;
        RECT  9.590 2.750 11.930 2.990 ;
        RECT  14.030 1.970 14.270 3.210 ;
        RECT  11.230 2.970 14.270 3.210 ;
        RECT  11.230 2.750 11.470 4.360 ;
        RECT  15.520 1.410 16.100 1.650 ;
        RECT  15.520 1.410 15.760 3.010 ;
        RECT  15.040 1.330 15.280 2.530 ;
        RECT  14.770 2.290 15.280 2.530 ;
        RECT  14.770 2.290 15.020 3.490 ;
        RECT  16.870 2.070 17.110 3.490 ;
        RECT  14.770 3.250 17.110 3.490 ;
        RECT  17.180 1.330 17.600 1.800 ;
        RECT  16.340 1.560 17.600 1.800 ;
        RECT  16.340 1.560 16.580 2.180 ;
        RECT  16.000 1.940 16.580 2.180 ;
        RECT  17.360 2.120 18.230 2.520 ;
        RECT  17.360 1.330 17.600 3.970 ;
        RECT  16.930 3.730 17.600 3.970 ;
    END
END slclq2

MACRO slclq1
    CLASS CORE ;
    FOREIGN slclq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.070 2.020 10.540 2.510 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.190 2.280 5.370 2.520 ;
        RECT  5.130 1.160 5.370 2.520 ;
        RECT  4.410 1.160 5.370 1.400 ;
        RECT  3.100 0.980 4.650 1.220 ;
        RECT  4.190 2.280 4.430 3.170 ;
        RECT  3.980 2.580 4.430 3.170 ;
        RECT  3.690 2.930 4.090 3.490 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.404  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 2.530 6.420 3.020 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.069  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.570 1.080 13.080 1.500 ;
        RECT  12.220 1.460 12.820 1.900 ;
        RECT  12.220 2.490 12.810 2.730 ;
        RECT  12.220 1.460 12.460 2.730 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.320 2.300 0.720 2.700 ;
        RECT  0.120 2.460 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.580 3.330 3.320 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.652  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.880 1.020 18.280 4.010 ;
        RECT  17.420 1.460 18.280 1.930 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 18.480 5.600 ;
        RECT  17.080 4.620 17.480 5.600 ;
        RECT  15.450 4.000 15.690 5.600 ;
        RECT  13.220 4.780 13.750 5.600 ;
        RECT  12.240 3.450 12.480 5.600 ;
        RECT  11.810 3.450 12.480 3.690 ;
        RECT  9.870 3.880 10.110 5.600 ;
        RECT  6.530 4.710 6.930 5.600 ;
        RECT  4.440 4.620 4.840 5.600 ;
        RECT  2.080 4.450 2.320 5.600 ;
        RECT  0.730 4.580 1.130 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 18.480 0.740 ;
        RECT  17.220 0.000 17.460 1.150 ;
        RECT  15.780 0.000 16.020 1.320 ;
        RECT  13.750 0.000 14.270 0.820 ;
        RECT  12.020 0.000 12.260 1.210 ;
        RECT  10.490 1.060 11.040 1.300 ;
        RECT  10.800 0.000 11.040 1.300 ;
        RECT  6.340 0.000 6.740 0.890 ;
        RECT  5.250 0.000 5.650 0.890 ;
        RECT  0.690 0.000 0.930 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.200 1.820 ;
        RECT  0.960 2.410 1.490 2.810 ;
        RECT  0.960 1.580 1.200 3.500 ;
        RECT  0.150 3.260 1.200 3.500 ;
        RECT  0.150 3.260 0.560 3.660 ;
        RECT  1.510 1.530 2.020 1.930 ;
        RECT  1.750 1.530 2.020 4.160 ;
        RECT  1.780 0.980 2.020 4.160 ;
        RECT  1.470 3.760 2.020 4.160 ;
        RECT  2.260 0.980 2.860 1.220 ;
        RECT  2.620 0.980 2.860 1.700 ;
        RECT  2.620 1.460 4.160 1.700 ;
        RECT  3.920 1.640 4.890 1.880 ;
        RECT  4.480 1.640 4.890 2.040 ;
        RECT  5.750 1.850 6.530 2.090 ;
        RECT  6.290 2.050 7.020 2.290 ;
        RECT  6.780 2.050 7.020 3.540 ;
        RECT  5.880 3.300 7.020 3.540 ;
        RECT  7.260 0.980 8.020 1.220 ;
        RECT  7.110 1.390 7.510 1.800 ;
        RECT  7.260 2.580 7.860 2.980 ;
        RECT  7.260 0.980 7.510 3.620 ;
        RECT  7.810 1.470 8.390 1.870 ;
        RECT  2.330 1.940 3.680 2.180 ;
        RECT  8.150 1.470 8.390 3.630 ;
        RECT  7.880 3.220 8.390 3.630 ;
        RECT  2.330 1.940 2.570 4.020 ;
        RECT  2.330 3.780 5.580 4.020 ;
        RECT  7.880 3.220 8.120 4.100 ;
        RECT  5.180 3.860 8.120 4.100 ;
        RECT  5.180 3.780 5.580 4.450 ;
        RECT  9.110 1.470 9.690 1.710 ;
        RECT  9.110 1.470 9.350 3.630 ;
        RECT  9.110 3.230 10.930 3.630 ;
        RECT  8.630 0.980 10.190 1.220 ;
        RECT  9.950 0.980 10.190 1.780 ;
        RECT  9.950 1.540 11.030 1.780 ;
        RECT  10.790 1.540 11.030 2.430 ;
        RECT  10.790 2.190 11.450 2.430 ;
        RECT  8.630 0.980 8.870 4.310 ;
        RECT  8.450 3.900 8.870 4.310 ;
        RECT  11.280 0.980 11.520 1.950 ;
        RECT  11.280 1.710 11.930 1.950 ;
        RECT  13.560 1.330 13.800 2.210 ;
        RECT  13.290 1.970 13.800 2.210 ;
        RECT  9.590 2.150 9.830 2.990 ;
        RECT  11.690 1.710 11.930 3.210 ;
        RECT  9.590 2.750 11.930 2.990 ;
        RECT  13.290 1.970 13.530 3.210 ;
        RECT  11.230 2.970 13.530 3.210 ;
        RECT  11.230 2.750 11.470 4.360 ;
        RECT  14.780 1.410 15.360 1.650 ;
        RECT  14.780 1.410 15.020 3.010 ;
        RECT  14.300 1.330 14.540 2.530 ;
        RECT  14.030 2.290 14.540 2.530 ;
        RECT  14.030 2.290 14.280 3.490 ;
        RECT  16.130 2.070 16.370 3.490 ;
        RECT  14.030 3.250 16.370 3.490 ;
        RECT  16.440 1.330 16.860 1.800 ;
        RECT  15.600 1.560 16.860 1.800 ;
        RECT  15.600 1.560 15.840 2.180 ;
        RECT  15.260 1.940 15.840 2.180 ;
        RECT  16.620 2.450 17.490 2.850 ;
        RECT  16.620 1.330 16.860 3.970 ;
        RECT  16.190 3.730 16.860 3.970 ;
    END
END slclq1

MACRO slchq4
    CLASS CORE ;
    FOREIGN slchq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.140 2.020 10.620 2.460 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.190 2.280 5.360 2.520 ;
        RECT  5.120 1.160 5.360 2.520 ;
        RECT  4.410 1.160 5.360 1.400 ;
        RECT  3.130 0.980 4.650 1.220 ;
        RECT  4.190 2.280 4.430 3.170 ;
        RECT  3.990 2.580 4.430 3.170 ;
        RECT  3.690 2.930 4.090 3.410 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.404  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 2.530 6.420 3.020 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.676  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.160 3.050 14.490 3.290 ;
        RECT  14.250 1.100 14.490 3.290 ;
        RECT  13.160 2.490 13.400 3.290 ;
        RECT  12.250 2.490 13.400 2.730 ;
        RECT  12.250 1.460 13.010 1.900 ;
        RECT  12.770 1.100 13.010 1.900 ;
        RECT  12.250 1.460 12.490 2.730 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.720 2.700 ;
        RECT  0.120 2.300 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.580 3.330 3.320 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.759  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.160 3.880 21.550 4.120 ;
        RECT  21.310 1.090 21.550 4.120 ;
        RECT  19.600 1.460 20.150 1.930 ;
        RECT  19.830 1.020 20.070 1.930 ;
        RECT  19.600 1.460 19.840 4.120 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 21.840 5.600 ;
        RECT  21.210 4.620 21.610 5.600 ;
        RECT  19.900 4.620 20.300 5.600 ;
        RECT  18.590 4.620 18.990 5.600 ;
        RECT  17.320 3.790 17.560 5.600 ;
        RECT  14.570 4.200 14.810 5.600 ;
        RECT  13.450 4.040 13.690 5.600 ;
        RECT  13.140 4.040 13.690 4.280 ;
        RECT  12.110 3.450 12.350 5.600 ;
        RECT  11.800 3.450 12.350 3.690 ;
        RECT  9.870 3.880 10.110 5.600 ;
        RECT  6.610 4.310 6.850 5.600 ;
        RECT  4.440 4.620 4.840 5.600 ;
        RECT  2.000 4.620 2.400 5.600 ;
        RECT  0.730 4.580 1.130 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 21.840 0.740 ;
        RECT  20.570 0.000 20.810 1.240 ;
        RECT  19.090 0.000 19.330 1.150 ;
        RECT  17.570 0.000 17.970 0.980 ;
        RECT  13.510 0.000 13.750 1.250 ;
        RECT  12.030 0.000 12.270 1.090 ;
        RECT  10.520 0.000 10.920 0.890 ;
        RECT  7.150 0.000 7.550 0.820 ;
        RECT  6.340 0.000 6.740 0.890 ;
        RECT  5.250 0.000 5.650 0.890 ;
        RECT  0.690 0.000 0.930 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.200 1.820 ;
        RECT  0.960 2.410 1.490 2.820 ;
        RECT  0.960 1.580 1.200 3.580 ;
        RECT  0.160 3.340 1.200 3.580 ;
        RECT  1.510 0.980 2.100 1.220 ;
        RECT  1.510 0.980 1.750 2.170 ;
        RECT  1.510 1.770 2.110 2.170 ;
        RECT  1.870 1.770 2.110 3.520 ;
        RECT  1.470 3.280 2.110 3.520 ;
        RECT  2.340 0.980 2.890 1.220 ;
        RECT  2.650 0.980 2.890 1.700 ;
        RECT  2.650 1.460 4.160 1.700 ;
        RECT  3.920 1.460 4.160 1.960 ;
        RECT  3.920 1.720 4.880 1.960 ;
        RECT  5.750 1.720 6.530 1.960 ;
        RECT  6.290 1.720 6.530 2.280 ;
        RECT  6.290 2.040 7.020 2.280 ;
        RECT  6.780 2.040 7.020 3.540 ;
        RECT  5.880 3.300 7.020 3.540 ;
        RECT  7.110 1.400 7.510 1.800 ;
        RECT  7.260 1.400 7.510 2.710 ;
        RECT  7.260 2.310 7.780 2.710 ;
        RECT  7.260 1.400 7.500 3.530 ;
        RECT  7.810 1.380 8.280 1.780 ;
        RECT  2.360 1.940 3.680 2.180 ;
        RECT  8.040 1.380 8.280 3.620 ;
        RECT  2.360 1.940 2.600 4.020 ;
        RECT  7.880 3.220 8.120 4.020 ;
        RECT  2.360 3.780 8.120 4.020 ;
        RECT  5.260 3.780 5.500 4.450 ;
        RECT  9.110 1.460 9.690 1.700 ;
        RECT  9.110 1.460 9.350 2.770 ;
        RECT  9.040 2.530 9.280 3.550 ;
        RECT  9.040 3.310 10.930 3.550 ;
        RECT  8.630 0.980 10.170 1.220 ;
        RECT  9.930 0.980 10.170 1.780 ;
        RECT  9.930 1.540 11.100 1.780 ;
        RECT  8.630 0.980 8.870 2.080 ;
        RECT  10.860 1.540 11.100 2.410 ;
        RECT  10.860 2.170 11.440 2.410 ;
        RECT  8.530 1.840 8.770 4.300 ;
        RECT  11.210 1.070 11.770 1.310 ;
        RECT  15.430 0.990 15.670 1.870 ;
        RECT  15.160 1.630 15.670 1.870 ;
        RECT  11.530 1.070 11.770 1.930 ;
        RECT  9.590 2.150 9.830 3.070 ;
        RECT  11.680 1.690 11.920 3.210 ;
        RECT  9.590 2.830 11.920 3.070 ;
        RECT  11.220 2.970 12.860 3.210 ;
        RECT  12.620 2.970 12.860 3.800 ;
        RECT  15.160 1.630 15.400 3.800 ;
        RECT  12.620 3.560 15.400 3.800 ;
        RECT  11.220 2.830 11.460 4.360 ;
        RECT  16.650 1.070 17.230 1.310 ;
        RECT  16.650 1.070 16.890 2.570 ;
        RECT  16.640 2.330 16.880 2.960 ;
        RECT  16.170 0.990 16.410 2.190 ;
        RECT  15.900 1.950 16.410 2.190 ;
        RECT  17.360 2.080 18.220 2.320 ;
        RECT  15.900 1.950 16.140 3.440 ;
        RECT  17.360 2.080 17.600 3.440 ;
        RECT  15.900 3.200 17.600 3.440 ;
        RECT  18.390 0.990 18.630 1.840 ;
        RECT  17.130 1.600 18.730 1.840 ;
        RECT  18.490 2.200 19.360 2.440 ;
        RECT  18.490 1.600 18.730 2.850 ;
        RECT  17.890 2.610 18.730 2.850 ;
    END
END slchq4

MACRO slchq2
    CLASS CORE ;
    FOREIGN slchq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.140 2.020 10.620 2.460 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.190 2.280 5.360 2.520 ;
        RECT  5.120 1.160 5.360 2.520 ;
        RECT  4.410 1.160 5.360 1.400 ;
        RECT  3.130 0.980 4.650 1.220 ;
        RECT  4.190 2.280 4.430 3.170 ;
        RECT  3.980 2.580 4.430 3.170 ;
        RECT  3.690 2.930 4.090 3.410 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.404  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 2.530 6.420 3.020 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.336  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.250 1.460 13.000 1.900 ;
        RECT  12.760 0.980 13.000 1.900 ;
        RECT  12.250 2.490 12.800 2.730 ;
        RECT  12.250 1.460 12.490 2.730 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.720 2.700 ;
        RECT  0.120 2.300 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.580 3.330 3.320 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.542  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.540 1.450 18.910 1.900 ;
        RECT  18.000 2.790 18.810 3.040 ;
        RECT  18.570 1.450 18.810 3.040 ;
        RECT  18.000 2.790 18.240 4.350 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.040 5.600 ;
        RECT  18.570 3.280 18.810 5.600 ;
        RECT  17.350 4.620 17.750 5.600 ;
        RECT  16.000 4.620 16.400 5.600 ;
        RECT  13.210 3.910 13.450 5.600 ;
        RECT  12.110 3.450 12.350 5.600 ;
        RECT  11.800 3.450 12.350 3.690 ;
        RECT  9.870 3.880 10.110 5.600 ;
        RECT  6.610 4.310 6.850 5.600 ;
        RECT  4.440 4.620 4.840 5.600 ;
        RECT  2.000 4.620 2.400 5.600 ;
        RECT  0.730 4.580 1.130 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.040 0.740 ;
        RECT  17.750 0.000 18.150 0.980 ;
        RECT  16.470 0.000 16.870 0.890 ;
        RECT  13.500 0.000 13.740 1.110 ;
        RECT  12.020 0.000 12.260 1.110 ;
        RECT  10.520 0.000 10.920 0.890 ;
        RECT  7.150 0.000 7.550 0.820 ;
        RECT  6.340 0.000 6.740 0.890 ;
        RECT  5.250 0.000 5.650 0.890 ;
        RECT  0.690 0.000 0.930 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.200 1.820 ;
        RECT  0.960 2.410 1.490 2.820 ;
        RECT  0.960 1.580 1.200 3.580 ;
        RECT  0.160 3.340 1.200 3.580 ;
        RECT  1.510 0.980 2.100 1.220 ;
        RECT  1.510 0.980 1.750 2.170 ;
        RECT  1.510 1.770 2.110 2.170 ;
        RECT  1.870 1.770 2.110 3.520 ;
        RECT  1.470 3.280 2.110 3.520 ;
        RECT  2.340 0.980 2.890 1.220 ;
        RECT  2.650 0.980 2.890 1.700 ;
        RECT  2.650 1.460 4.160 1.700 ;
        RECT  3.920 1.460 4.160 1.960 ;
        RECT  3.920 1.720 4.880 1.960 ;
        RECT  5.750 1.720 6.530 1.960 ;
        RECT  6.290 1.720 6.530 2.280 ;
        RECT  6.290 2.040 7.020 2.280 ;
        RECT  6.780 2.040 7.020 3.540 ;
        RECT  5.880 3.300 7.020 3.540 ;
        RECT  7.110 1.400 7.510 1.800 ;
        RECT  7.260 1.400 7.510 2.710 ;
        RECT  7.260 2.310 7.780 2.710 ;
        RECT  7.260 1.400 7.500 3.530 ;
        RECT  7.810 1.380 8.280 1.780 ;
        RECT  2.360 1.940 3.680 2.180 ;
        RECT  8.040 1.380 8.280 3.620 ;
        RECT  2.360 1.940 2.600 4.020 ;
        RECT  7.880 3.220 8.120 4.020 ;
        RECT  2.360 3.780 8.120 4.020 ;
        RECT  5.260 3.780 5.500 4.450 ;
        RECT  9.110 1.460 9.690 1.700 ;
        RECT  9.110 1.460 9.350 2.770 ;
        RECT  9.040 2.530 9.280 3.550 ;
        RECT  9.040 3.310 10.930 3.550 ;
        RECT  8.630 0.980 10.170 1.220 ;
        RECT  9.930 0.980 10.170 1.780 ;
        RECT  9.930 1.540 11.100 1.780 ;
        RECT  8.630 0.980 8.870 2.080 ;
        RECT  10.860 1.540 11.100 2.410 ;
        RECT  10.860 2.170 11.440 2.410 ;
        RECT  8.530 1.840 8.770 4.300 ;
        RECT  11.200 1.070 11.770 1.310 ;
        RECT  14.300 1.100 14.540 1.670 ;
        RECT  13.920 1.430 14.540 1.670 ;
        RECT  11.530 1.070 11.770 1.930 ;
        RECT  9.590 2.150 9.830 3.070 ;
        RECT  11.680 1.690 11.920 3.210 ;
        RECT  9.590 2.830 11.920 3.070 ;
        RECT  11.220 2.970 14.160 3.210 ;
        RECT  13.920 1.430 14.160 3.630 ;
        RECT  11.220 2.830 11.460 4.360 ;
        RECT  15.780 1.100 16.020 2.020 ;
        RECT  15.280 1.780 16.020 2.020 ;
        RECT  15.280 1.780 15.520 3.090 ;
        RECT  15.400 2.850 15.640 3.630 ;
        RECT  14.780 1.100 15.360 1.500 ;
        RECT  14.780 1.100 15.020 2.150 ;
        RECT  16.120 2.780 16.880 3.020 ;
        RECT  14.660 1.910 14.900 4.130 ;
        RECT  16.120 2.780 16.360 4.130 ;
        RECT  14.660 3.880 16.360 4.130 ;
        RECT  15.790 2.300 17.360 2.540 ;
        RECT  17.120 1.770 17.360 2.540 ;
        RECT  17.250 2.310 18.220 2.550 ;
        RECT  17.250 2.310 17.490 3.550 ;
        RECT  16.650 3.310 17.490 3.550 ;
    END
END slchq2

MACRO slchq1
    CLASS CORE ;
    FOREIGN slchq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.140 2.020 10.620 2.460 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.190 2.280 5.360 2.520 ;
        RECT  5.120 1.160 5.360 2.520 ;
        RECT  4.410 1.160 5.360 1.400 ;
        RECT  3.130 0.980 4.650 1.220 ;
        RECT  4.190 2.280 4.430 3.170 ;
        RECT  3.980 2.580 4.430 3.170 ;
        RECT  3.690 2.930 4.090 3.410 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.404  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 2.530 6.420 3.020 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.069  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.250 1.460 13.000 1.900 ;
        RECT  12.760 0.980 13.000 1.900 ;
        RECT  12.250 2.490 12.800 2.730 ;
        RECT  12.250 1.460 12.490 2.730 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.720 2.700 ;
        RECT  0.120 2.300 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.580 3.330 3.320 ;
        END
    END SD
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.340 3.080 17.800 3.580 ;
        RECT  17.560 1.310 17.800 3.580 ;
        RECT  17.100 1.310 17.800 1.550 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.920 5.600 ;
        RECT  16.770 4.620 17.170 5.600 ;
        RECT  15.420 4.620 15.820 5.600 ;
        RECT  12.110 3.450 12.350 5.600 ;
        RECT  11.800 3.450 12.350 3.690 ;
        RECT  9.870 3.880 10.110 5.600 ;
        RECT  6.610 4.310 6.850 5.600 ;
        RECT  4.440 4.620 4.840 5.600 ;
        RECT  2.000 4.620 2.400 5.600 ;
        RECT  0.730 4.580 1.130 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.920 0.740 ;
        RECT  16.970 0.000 17.370 0.890 ;
        RECT  15.740 0.000 16.140 0.890 ;
        RECT  12.020 0.000 12.260 1.110 ;
        RECT  10.520 0.000 10.920 0.890 ;
        RECT  7.150 0.000 7.550 0.820 ;
        RECT  6.340 0.000 6.740 0.890 ;
        RECT  5.250 0.000 5.650 0.890 ;
        RECT  0.690 0.000 0.930 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.200 1.820 ;
        RECT  0.960 2.410 1.490 2.820 ;
        RECT  0.960 1.580 1.200 3.580 ;
        RECT  0.160 3.340 1.200 3.580 ;
        RECT  1.510 0.980 2.100 1.220 ;
        RECT  1.510 0.980 1.750 2.170 ;
        RECT  1.510 1.770 2.110 2.170 ;
        RECT  1.870 1.770 2.110 3.520 ;
        RECT  1.470 3.280 2.110 3.520 ;
        RECT  2.340 0.980 2.890 1.220 ;
        RECT  2.650 0.980 2.890 1.700 ;
        RECT  2.650 1.460 4.160 1.700 ;
        RECT  3.920 1.460 4.160 1.960 ;
        RECT  3.920 1.720 4.880 1.960 ;
        RECT  5.750 1.720 6.530 1.960 ;
        RECT  6.290 1.720 6.530 2.280 ;
        RECT  6.290 2.040 7.020 2.280 ;
        RECT  6.780 2.040 7.020 3.540 ;
        RECT  5.880 3.300 7.020 3.540 ;
        RECT  7.110 1.400 7.510 1.800 ;
        RECT  7.260 1.400 7.510 2.710 ;
        RECT  7.260 2.310 7.780 2.710 ;
        RECT  7.260 1.400 7.500 3.530 ;
        RECT  7.810 1.380 8.280 1.780 ;
        RECT  2.360 1.940 3.680 2.180 ;
        RECT  8.040 1.380 8.280 3.620 ;
        RECT  2.360 1.940 2.600 4.020 ;
        RECT  7.880 3.220 8.120 4.020 ;
        RECT  2.360 3.780 8.120 4.020 ;
        RECT  5.260 3.780 5.500 4.450 ;
        RECT  9.110 1.460 9.690 1.700 ;
        RECT  9.110 1.460 9.350 2.770 ;
        RECT  9.040 2.530 9.280 3.550 ;
        RECT  9.040 3.310 10.930 3.550 ;
        RECT  8.630 0.980 10.170 1.220 ;
        RECT  9.930 0.980 10.170 1.780 ;
        RECT  9.930 1.540 11.100 1.780 ;
        RECT  8.630 0.980 8.870 2.080 ;
        RECT  10.860 1.540 11.100 2.410 ;
        RECT  10.860 2.170 11.440 2.410 ;
        RECT  8.530 1.840 8.770 4.300 ;
        RECT  11.200 1.070 11.770 1.310 ;
        RECT  13.560 1.100 13.800 1.670 ;
        RECT  11.530 1.070 11.770 1.930 ;
        RECT  9.590 2.150 9.830 3.070 ;
        RECT  11.680 1.690 11.920 3.210 ;
        RECT  9.590 2.830 11.920 3.070 ;
        RECT  11.220 2.970 13.580 3.210 ;
        RECT  13.340 1.430 13.580 3.630 ;
        RECT  11.220 2.830 11.460 4.360 ;
        RECT  15.040 1.100 15.280 2.020 ;
        RECT  14.700 1.780 15.280 2.020 ;
        RECT  14.700 1.780 14.940 3.090 ;
        RECT  14.820 2.850 15.060 3.630 ;
        RECT  14.080 1.100 14.620 1.500 ;
        RECT  15.540 2.780 16.300 3.020 ;
        RECT  14.080 1.100 14.320 4.130 ;
        RECT  15.540 2.780 15.780 4.130 ;
        RECT  14.080 3.880 15.780 4.130 ;
        RECT  16.380 1.770 16.620 2.540 ;
        RECT  15.210 2.300 16.910 2.540 ;
        RECT  16.670 2.580 17.320 2.840 ;
        RECT  16.670 2.300 16.910 3.550 ;
        RECT  16.070 3.310 16.910 3.550 ;
    END
END slchq1

MACRO slbhb4
    CLASS CORE ;
    FOREIGN slbhb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 28.560 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.477  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.350 2.740 3.020 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.390 2.020 5.630 2.770 ;
        RECT  5.100 2.020 5.630 2.460 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.404  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  27.870 2.930 28.440 3.330 ;
        RECT  28.060 2.330 28.440 3.330 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.756  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.290 3.140 18.980 3.580 ;
        RECT  16.910 2.960 18.840 3.200 ;
        RECT  18.600 1.430 18.840 3.580 ;
        RECT  17.120 1.800 18.840 2.040 ;
        RECT  17.120 1.320 17.360 2.040 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.836  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.180 3.110 12.820 3.510 ;
        RECT  12.580 1.800 12.820 3.510 ;
        RECT  12.380 2.580 12.820 3.510 ;
        RECT  10.810 1.800 12.820 2.040 ;
        RECT  12.290 1.430 12.530 2.040 ;
        RECT  10.870 3.190 12.820 3.430 ;
        RECT  10.810 1.430 11.050 2.040 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.477  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.710 3.020 ;
        RECT  0.120 2.130 0.410 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.120 2.460 3.860 3.020 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.486  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.560 2.420 15.060 3.020 ;
        END
    END SDN
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.017  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  25.510 2.580 25.770 3.890 ;
        RECT  25.530 1.610 25.770 3.890 ;
        RECT  24.090 1.930 25.770 2.170 ;
        RECT  24.050 3.200 25.770 3.440 ;
        RECT  25.260 2.580 25.770 3.440 ;
        RECT  24.090 1.700 24.490 2.170 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 28.560 5.600 ;
        RECT  27.440 4.540 27.840 5.600 ;
        RECT  26.170 4.620 26.570 5.600 ;
        RECT  24.870 4.620 25.270 5.600 ;
        RECT  23.480 4.610 23.880 5.600 ;
        RECT  22.000 4.640 22.400 5.600 ;
        RECT  19.060 4.710 19.460 5.600 ;
        RECT  17.700 4.710 18.100 5.600 ;
        RECT  16.220 4.710 16.620 5.600 ;
        RECT  14.920 4.710 15.320 5.600 ;
        RECT  13.560 4.710 13.960 5.600 ;
        RECT  12.780 4.710 13.180 5.600 ;
        RECT  11.420 4.710 11.830 5.600 ;
        RECT  9.920 4.710 10.320 5.600 ;
        RECT  7.760 4.710 8.160 5.600 ;
        RECT  4.250 4.400 4.490 5.600 ;
        RECT  2.280 4.400 2.520 5.600 ;
        RECT  0.800 4.160 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 28.560 0.740 ;
        RECT  27.720 0.000 27.960 1.180 ;
        RECT  24.860 0.000 25.260 0.890 ;
        RECT  23.270 0.000 23.670 0.890 ;
        RECT  22.610 0.000 23.010 0.890 ;
        RECT  19.340 0.000 19.580 1.640 ;
        RECT  17.620 1.320 18.180 1.560 ;
        RECT  17.620 0.000 17.860 1.560 ;
        RECT  16.370 0.000 16.610 1.640 ;
        RECT  14.930 0.000 15.170 1.640 ;
        RECT  12.790 1.320 13.350 1.560 ;
        RECT  12.790 0.000 13.030 1.560 ;
        RECT  11.320 1.310 11.870 1.560 ;
        RECT  11.320 0.000 11.560 1.560 ;
        RECT  10.070 0.000 10.310 1.640 ;
        RECT  8.630 0.000 8.870 1.670 ;
        RECT  2.030 0.000 2.430 0.890 ;
        RECT  0.730 0.000 1.130 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.210 1.820 ;
        RECT  0.970 2.110 1.530 2.350 ;
        RECT  0.970 1.580 1.210 3.520 ;
        RECT  0.150 3.280 1.210 3.520 ;
        RECT  2.800 0.980 4.940 1.220 ;
        RECT  2.800 0.980 3.200 1.410 ;
        RECT  1.510 1.230 2.010 1.630 ;
        RECT  1.770 1.870 3.390 2.110 ;
        RECT  1.770 1.230 2.010 2.940 ;
        RECT  4.100 2.760 5.030 3.000 ;
        RECT  4.100 2.760 4.340 3.500 ;
        RECT  1.480 3.260 4.340 3.500 ;
        RECT  1.480 2.620 1.900 3.580 ;
        RECT  5.840 1.020 6.080 1.700 ;
        RECT  4.110 1.460 6.110 1.700 ;
        RECT  4.110 1.460 4.350 2.120 ;
        RECT  5.870 1.460 6.110 3.470 ;
        RECT  5.270 3.070 6.110 3.470 ;
        RECT  5.270 3.070 5.510 4.050 ;
        RECT  2.770 3.810 5.510 4.050 ;
        RECT  7.310 2.180 7.550 2.980 ;
        RECT  7.310 2.740 8.980 2.980 ;
        RECT  7.350 1.330 7.590 1.880 ;
        RECT  6.830 1.640 8.390 1.880 ;
        RECT  8.150 1.640 8.390 2.310 ;
        RECT  8.150 2.070 9.350 2.310 ;
        RECT  9.110 2.310 9.490 2.510 ;
        RECT  9.160 2.470 9.810 2.540 ;
        RECT  9.220 2.470 9.810 2.710 ;
        RECT  6.830 1.640 7.070 3.510 ;
        RECT  6.830 3.270 9.020 3.510 ;
        RECT  9.250 1.620 9.830 1.830 ;
        RECT  9.250 1.590 9.710 1.830 ;
        RECT  9.590 1.810 9.900 2.050 ;
        RECT  9.690 1.930 10.290 2.170 ;
        RECT  10.050 2.300 11.990 2.700 ;
        RECT  10.050 1.930 10.290 3.260 ;
        RECT  9.330 3.020 10.290 3.260 ;
        RECT  6.350 1.130 6.910 1.370 ;
        RECT  13.870 2.410 14.270 2.940 ;
        RECT  13.850 2.700 14.090 3.990 ;
        RECT  6.160 3.750 14.090 3.990 ;
        RECT  6.350 1.130 6.590 4.140 ;
        RECT  6.160 3.740 6.590 4.140 ;
        RECT  13.650 1.320 14.610 1.580 ;
        RECT  14.370 1.320 14.610 2.120 ;
        RECT  14.370 1.880 15.540 2.120 ;
        RECT  15.300 2.340 15.850 2.580 ;
        RECT  15.300 1.880 15.540 3.500 ;
        RECT  14.330 3.260 15.540 3.500 ;
        RECT  15.550 1.240 16.130 1.640 ;
        RECT  15.830 1.820 16.190 2.100 ;
        RECT  15.830 1.240 16.130 2.100 ;
        RECT  16.090 2.280 16.960 2.680 ;
        RECT  16.090 1.880 16.330 3.990 ;
        RECT  15.620 3.750 16.330 3.990 ;
        RECT  19.660 2.260 20.290 2.500 ;
        RECT  20.040 1.450 20.290 3.650 ;
        RECT  19.860 3.250 20.290 3.650 ;
        RECT  21.350 1.460 21.840 1.860 ;
        RECT  21.350 1.460 21.590 2.500 ;
        RECT  21.100 2.260 21.590 2.500 ;
        RECT  21.100 2.260 21.340 3.410 ;
        RECT  21.100 3.170 21.830 3.410 ;
        RECT  20.550 1.590 21.100 1.830 ;
        RECT  22.600 2.590 22.840 3.250 ;
        RECT  22.070 3.010 22.840 3.250 ;
        RECT  20.550 1.590 20.790 4.100 ;
        RECT  22.070 3.010 22.310 3.890 ;
        RECT  20.550 3.650 22.310 3.890 ;
        RECT  20.550 3.650 21.050 4.100 ;
        RECT  22.470 1.610 23.350 1.850 ;
        RECT  22.470 1.610 22.710 2.330 ;
        RECT  21.910 2.090 22.710 2.330 ;
        RECT  21.910 2.090 22.150 2.770 ;
        RECT  23.110 2.410 24.900 2.810 ;
        RECT  23.110 1.610 23.350 3.730 ;
        RECT  22.770 3.490 23.350 3.730 ;
        RECT  26.510 1.000 26.770 1.620 ;
        RECT  26.730 1.380 26.970 2.540 ;
        RECT  26.490 2.300 26.730 3.810 ;
        RECT  26.490 3.570 27.100 3.810 ;
        RECT  20.450 0.980 22.300 1.220 ;
        RECT  22.070 1.130 26.250 1.370 ;
        RECT  27.390 1.840 28.410 2.080 ;
        RECT  27.070 3.040 27.630 3.280 ;
        RECT  27.390 3.610 28.410 3.850 ;
        RECT  26.010 1.130 26.250 4.370 ;
        RECT  26.600 4.050 27.630 4.290 ;
        RECT  22.720 4.130 27.630 4.290 ;
        RECT  27.390 1.840 27.630 4.290 ;
        RECT  21.330 4.150 26.840 4.370 ;
        RECT  21.330 4.150 22.960 4.390 ;
        RECT  7.190 4.230 20.250 4.470 ;
        RECT  5.930 4.380 7.420 4.620 ;
        RECT  20.020 4.380 21.570 4.620 ;
    END
END slbhb4

MACRO slbhb2
    CLASS CORE ;
    FOREIGN slbhb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.477  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.350 2.740 3.020 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.390 2.020 5.630 2.770 ;
        RECT  5.100 2.020 5.630 2.460 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  23.510 2.330 23.960 3.580 ;
        RECT  23.200 2.930 23.960 3.330 ;
        RECT  23.450 2.330 23.960 3.330 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.119  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.660 3.580 16.060 3.980 ;
        RECT  15.180 3.140 15.670 3.860 ;
        RECT  15.430 1.380 15.670 3.860 ;
        RECT  14.360 3.620 16.060 3.860 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.570  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.700 3.090 11.270 3.490 ;
        RECT  10.700 2.580 11.140 3.490 ;
        RECT  10.900 1.460 11.140 3.490 ;
        RECT  10.730 1.460 11.140 1.900 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.477  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.710 3.020 ;
        RECT  0.120 2.130 0.410 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.120 2.460 3.860 3.020 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.479  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.800 2.020 12.260 2.720 ;
        END
    END SDN
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.555  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  20.470 2.020 21.320 2.460 ;
        RECT  20.920 1.690 21.320 2.460 ;
        RECT  20.470 3.170 21.020 3.410 ;
        RECT  20.470 2.020 20.710 3.410 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 24.080 5.600 ;
        RECT  22.640 4.610 23.060 5.600 ;
        RECT  21.360 4.620 21.760 5.600 ;
        RECT  20.050 4.620 20.450 5.600 ;
        RECT  18.720 4.640 19.110 5.600 ;
        RECT  14.950 4.710 15.350 5.600 ;
        RECT  13.050 4.710 13.450 5.600 ;
        RECT  11.540 4.710 11.940 5.600 ;
        RECT  9.920 4.710 10.320 5.600 ;
        RECT  7.760 4.710 8.160 5.600 ;
        RECT  4.250 4.400 4.490 5.600 ;
        RECT  2.280 4.400 2.520 5.600 ;
        RECT  0.800 4.160 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 24.080 0.740 ;
        RECT  23.210 0.000 23.610 1.180 ;
        RECT  20.080 0.000 20.480 0.890 ;
        RECT  19.440 0.000 19.840 0.890 ;
        RECT  15.940 1.320 16.490 1.560 ;
        RECT  15.940 0.000 16.180 1.560 ;
        RECT  14.600 1.320 15.150 1.560 ;
        RECT  14.910 0.000 15.150 1.560 ;
        RECT  11.550 0.000 11.790 1.640 ;
        RECT  10.070 0.000 10.310 1.640 ;
        RECT  8.630 0.000 8.870 1.670 ;
        RECT  2.030 0.000 2.430 0.890 ;
        RECT  0.730 0.000 1.130 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.210 1.820 ;
        RECT  0.970 2.110 1.530 2.350 ;
        RECT  0.970 1.580 1.210 3.520 ;
        RECT  0.150 3.280 1.210 3.520 ;
        RECT  2.800 0.980 4.940 1.220 ;
        RECT  2.800 0.980 3.200 1.410 ;
        RECT  1.510 1.230 2.010 1.630 ;
        RECT  1.770 1.870 3.390 2.110 ;
        RECT  1.770 1.230 2.010 2.940 ;
        RECT  4.100 2.760 5.030 3.000 ;
        RECT  4.100 2.760 4.340 3.500 ;
        RECT  1.480 3.260 4.340 3.500 ;
        RECT  1.480 2.620 1.900 3.580 ;
        RECT  5.840 1.020 6.080 1.700 ;
        RECT  4.110 1.460 6.110 1.700 ;
        RECT  4.110 1.460 4.350 2.120 ;
        RECT  5.870 1.460 6.110 3.470 ;
        RECT  5.270 3.070 6.110 3.470 ;
        RECT  5.270 3.070 5.510 4.050 ;
        RECT  2.770 3.810 5.510 4.050 ;
        RECT  7.310 2.180 7.550 2.980 ;
        RECT  7.310 2.740 8.980 2.980 ;
        RECT  7.350 1.330 7.590 1.880 ;
        RECT  6.830 1.640 8.390 1.880 ;
        RECT  8.150 1.640 8.390 2.310 ;
        RECT  8.150 2.070 9.350 2.310 ;
        RECT  9.110 2.310 9.490 2.510 ;
        RECT  9.160 2.470 9.790 2.540 ;
        RECT  9.220 2.470 9.790 2.710 ;
        RECT  6.830 1.640 7.070 3.510 ;
        RECT  6.830 3.270 9.020 3.510 ;
        RECT  9.250 1.620 9.830 1.830 ;
        RECT  9.250 1.590 9.710 1.830 ;
        RECT  9.590 1.810 9.900 2.050 ;
        RECT  9.690 1.930 10.290 2.170 ;
        RECT  10.050 2.120 10.600 2.360 ;
        RECT  10.050 1.930 10.290 3.260 ;
        RECT  9.330 3.020 10.290 3.260 ;
        RECT  6.350 1.130 6.910 1.370 ;
        RECT  12.640 2.190 12.880 3.230 ;
        RECT  11.630 2.990 12.880 3.230 ;
        RECT  11.630 2.990 11.870 3.990 ;
        RECT  6.160 3.750 11.870 3.990 ;
        RECT  6.350 1.130 6.590 4.140 ;
        RECT  6.160 3.740 6.590 4.140 ;
        RECT  13.130 2.340 13.810 2.580 ;
        RECT  13.130 1.550 13.370 3.840 ;
        RECT  12.310 3.600 13.370 3.840 ;
        RECT  13.860 1.240 14.320 1.640 ;
        RECT  14.080 1.240 14.320 2.100 ;
        RECT  14.080 1.860 14.680 2.100 ;
        RECT  14.440 2.120 15.190 2.360 ;
        RECT  14.440 1.860 14.680 3.060 ;
        RECT  13.730 2.820 14.680 3.060 ;
        RECT  13.730 2.820 13.970 3.420 ;
        RECT  16.870 1.430 17.120 2.040 ;
        RECT  16.670 1.800 16.910 3.690 ;
        RECT  16.260 2.750 16.910 3.160 ;
        RECT  16.470 2.750 16.910 3.690 ;
        RECT  18.170 1.460 18.670 1.860 ;
        RECT  18.100 1.920 18.220 2.230 ;
        RECT  18.070 1.950 18.410 2.140 ;
        RECT  18.170 1.460 18.410 2.140 ;
        RECT  17.860 1.990 18.290 2.170 ;
        RECT  17.860 1.990 18.240 2.180 ;
        RECT  17.860 1.990 18.100 2.930 ;
        RECT  17.790 2.710 18.100 2.930 ;
        RECT  17.720 2.760 17.960 3.430 ;
        RECT  17.720 3.190 18.440 3.430 ;
        RECT  17.380 1.510 17.930 1.750 ;
        RECT  17.380 1.510 17.620 2.520 ;
        RECT  18.920 3.010 19.470 3.250 ;
        RECT  19.230 2.580 19.470 3.250 ;
        RECT  17.150 2.280 17.390 4.100 ;
        RECT  18.850 3.070 19.090 3.910 ;
        RECT  17.150 3.670 19.090 3.910 ;
        RECT  17.150 3.670 17.650 4.100 ;
        RECT  19.630 1.610 20.030 2.340 ;
        RECT  18.670 2.100 20.030 2.340 ;
        RECT  19.750 1.610 20.030 2.820 ;
        RECT  18.670 2.100 18.910 2.620 ;
        RECT  18.410 2.380 18.910 2.620 ;
        RECT  19.750 2.420 20.230 2.820 ;
        RECT  18.410 2.380 18.650 2.930 ;
        RECT  19.750 1.610 19.990 3.730 ;
        RECT  19.330 3.490 19.990 3.730 ;
        RECT  22.100 1.530 22.340 2.160 ;
        RECT  21.730 2.450 22.180 2.850 ;
        RECT  21.940 1.920 22.180 3.890 ;
        RECT  21.940 3.460 22.460 3.890 ;
        RECT  17.340 0.980 19.130 1.220 ;
        RECT  21.400 0.980 22.950 1.220 ;
        RECT  18.900 1.130 21.630 1.370 ;
        RECT  22.710 1.840 23.800 2.080 ;
        RECT  22.710 0.980 22.950 2.650 ;
        RECT  22.600 2.400 22.940 3.220 ;
        RECT  22.440 2.820 22.940 3.220 ;
        RECT  22.700 2.400 22.940 4.370 ;
        RECT  19.550 4.130 23.800 4.370 ;
        RECT  18.220 4.150 19.790 4.390 ;
        RECT  7.190 4.230 16.540 4.470 ;
        RECT  5.930 4.380 7.420 4.620 ;
        RECT  16.310 4.380 18.460 4.620 ;
    END
END slbhb2

MACRO slbhb1
    CLASS CORE ;
    FOREIGN slbhb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.477  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.350 2.740 3.020 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.390 2.020 5.630 2.770 ;
        RECT  5.100 2.020 5.630 2.460 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  21.900 2.930 22.280 3.580 ;
        RECT  21.920 2.330 22.280 3.580 ;
        RECT  21.550 2.930 22.280 3.330 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.222  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.020 1.720 15.260 2.910 ;
        RECT  14.940 1.380 15.180 1.900 ;
        RECT  14.620 3.130 15.150 3.580 ;
        RECT  14.750 2.660 15.150 3.580 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.224  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.700 3.090 11.270 3.490 ;
        RECT  10.700 2.580 11.140 3.490 ;
        RECT  10.900 1.460 11.140 3.490 ;
        RECT  10.730 1.460 11.140 1.900 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.477  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.710 3.020 ;
        RECT  0.120 2.130 0.410 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.120 2.460 3.860 3.020 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.380 2.420 12.820 3.020 ;
        END
    END SDN
    PIN SO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.120  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.520 1.700 20.100 2.460 ;
        RECT  19.520 3.660 20.070 3.900 ;
        RECT  19.520 1.700 19.760 3.900 ;
        END
    END SO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 22.400 5.600 ;
        RECT  20.980 4.620 21.380 5.600 ;
        RECT  19.100 4.620 19.500 5.600 ;
        RECT  17.620 4.710 18.020 5.600 ;
        RECT  14.040 4.710 14.440 5.600 ;
        RECT  12.740 4.710 13.140 5.600 ;
        RECT  11.220 4.710 11.620 5.600 ;
        RECT  9.920 4.710 10.320 5.600 ;
        RECT  7.760 4.710 8.160 5.600 ;
        RECT  4.250 4.400 4.490 5.600 ;
        RECT  2.280 4.400 2.520 5.600 ;
        RECT  0.800 4.160 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 22.400 0.740 ;
        RECT  21.600 0.000 22.010 0.890 ;
        RECT  18.300 0.000 18.700 0.890 ;
        RECT  14.110 1.320 14.680 1.560 ;
        RECT  14.440 0.000 14.680 1.560 ;
        RECT  12.740 0.000 13.000 1.640 ;
        RECT  10.070 0.000 10.310 1.640 ;
        RECT  8.630 0.000 8.870 1.670 ;
        RECT  2.030 0.000 2.430 0.890 ;
        RECT  0.730 0.000 1.130 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.210 1.820 ;
        RECT  0.970 2.110 1.530 2.350 ;
        RECT  0.970 1.580 1.210 3.520 ;
        RECT  0.150 3.280 1.210 3.520 ;
        RECT  2.800 0.980 4.940 1.220 ;
        RECT  2.800 0.980 3.200 1.410 ;
        RECT  1.510 1.230 2.010 1.630 ;
        RECT  1.770 1.870 3.390 2.110 ;
        RECT  1.770 1.230 2.010 2.940 ;
        RECT  4.100 2.760 5.030 3.000 ;
        RECT  4.100 2.760 4.340 3.500 ;
        RECT  1.480 3.260 4.340 3.500 ;
        RECT  1.480 2.620 1.900 3.580 ;
        RECT  5.840 1.020 6.080 1.700 ;
        RECT  4.110 1.460 6.110 1.700 ;
        RECT  4.110 1.460 4.350 2.120 ;
        RECT  5.870 1.460 6.110 3.460 ;
        RECT  5.270 3.060 6.110 3.460 ;
        RECT  5.270 3.060 5.510 4.050 ;
        RECT  2.770 3.810 5.510 4.050 ;
        RECT  7.310 2.180 7.550 2.980 ;
        RECT  7.310 2.740 8.980 2.980 ;
        RECT  7.350 1.330 7.590 1.880 ;
        RECT  6.830 1.640 8.390 1.880 ;
        RECT  8.150 1.640 8.390 2.310 ;
        RECT  8.150 2.070 9.350 2.310 ;
        RECT  9.110 2.310 9.480 2.510 ;
        RECT  9.160 2.470 9.790 2.540 ;
        RECT  9.220 2.470 9.790 2.710 ;
        RECT  6.830 1.640 7.070 3.510 ;
        RECT  6.830 3.270 9.020 3.510 ;
        RECT  9.250 1.620 9.830 1.830 ;
        RECT  9.250 1.590 9.710 1.830 ;
        RECT  9.590 1.810 9.900 2.050 ;
        RECT  9.690 1.930 10.290 2.170 ;
        RECT  10.050 2.120 10.600 2.360 ;
        RECT  10.050 1.930 10.290 3.260 ;
        RECT  9.330 3.020 10.290 3.260 ;
        RECT  6.350 1.130 6.910 1.370 ;
        RECT  11.690 2.410 12.090 2.940 ;
        RECT  11.670 2.700 11.910 3.990 ;
        RECT  6.160 3.750 11.910 3.990 ;
        RECT  6.350 1.130 6.590 4.140 ;
        RECT  6.160 3.740 6.590 4.140 ;
        RECT  11.470 1.320 12.430 1.580 ;
        RECT  12.190 1.320 12.430 2.120 ;
        RECT  12.190 1.880 13.300 2.120 ;
        RECT  13.060 2.340 13.620 2.580 ;
        RECT  13.060 1.880 13.300 3.500 ;
        RECT  12.150 3.260 13.300 3.500 ;
        RECT  13.370 1.240 13.830 1.640 ;
        RECT  13.590 1.240 13.830 2.100 ;
        RECT  13.590 1.860 14.150 2.100 ;
        RECT  13.910 2.140 14.780 2.380 ;
        RECT  13.910 1.860 14.150 3.990 ;
        RECT  13.440 3.750 14.150 3.990 ;
        RECT  15.460 3.250 15.890 3.650 ;
        RECT  15.620 3.250 15.890 4.140 ;
        RECT  15.640 1.450 15.890 4.140 ;
        RECT  15.290 3.890 15.890 4.140 ;
        RECT  16.950 1.460 17.440 1.860 ;
        RECT  16.950 1.460 17.190 2.500 ;
        RECT  16.700 2.260 17.190 2.500 ;
        RECT  16.700 2.260 16.940 3.440 ;
        RECT  16.700 3.200 17.430 3.440 ;
        RECT  16.150 1.590 16.700 1.830 ;
        RECT  18.200 2.590 18.440 3.250 ;
        RECT  17.670 3.010 18.440 3.250 ;
        RECT  16.150 1.590 16.390 4.100 ;
        RECT  17.670 3.010 17.910 3.990 ;
        RECT  16.150 3.750 17.910 3.990 ;
        RECT  16.150 3.700 16.650 4.100 ;
        RECT  18.070 1.610 18.950 1.850 ;
        RECT  18.070 1.610 18.310 2.330 ;
        RECT  17.510 2.090 18.310 2.330 ;
        RECT  18.710 2.360 19.260 2.600 ;
        RECT  17.510 2.090 17.750 2.770 ;
        RECT  18.710 1.610 18.950 3.730 ;
        RECT  18.380 3.490 18.950 3.730 ;
        RECT  20.490 1.530 20.890 2.160 ;
        RECT  20.150 2.750 20.580 3.150 ;
        RECT  20.340 3.370 20.670 3.580 ;
        RECT  20.340 1.920 20.580 3.580 ;
        RECT  20.380 3.460 20.780 3.890 ;
        RECT  16.050 0.980 18.070 1.220 ;
        RECT  18.950 0.980 21.370 1.220 ;
        RECT  17.840 1.130 19.180 1.370 ;
        RECT  21.130 1.840 22.250 2.080 ;
        RECT  21.130 0.980 21.370 2.650 ;
        RECT  20.860 2.820 21.260 3.220 ;
        RECT  21.020 2.400 21.260 4.380 ;
        RECT  7.190 4.230 14.900 4.470 ;
        RECT  17.110 4.230 22.200 4.380 ;
        RECT  18.150 4.140 22.200 4.380 ;
        RECT  5.930 4.380 18.390 4.470 ;
        RECT  5.930 4.380 7.420 4.620 ;
        RECT  14.670 4.380 17.350 4.620 ;
    END
END slbhb1

MACRO skbrb4
    CLASS CORE ;
    FOREIGN skbrb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 29.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.110 2.520 14.660 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.243  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 2.580 9.350 3.160 ;
        END
    END CP
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.369  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 5.070 2.480 ;
        END
    END J
    PIN KZ
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.020 7.740 2.600 ;
        END
    END KZ
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.574  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  27.680 2.580 28.140 4.180 ;
        RECT  27.740 1.770 28.140 4.180 ;
        RECT  26.380 2.580 28.140 3.020 ;
        RECT  26.380 1.770 26.780 4.150 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.619  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  24.960 2.530 25.420 4.180 ;
        RECT  25.020 1.770 25.420 4.180 ;
        RECT  23.570 2.530 25.420 3.020 ;
        RECT  23.660 1.770 24.060 4.150 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.340 0.700 2.740 ;
        RECT  0.120 2.340 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.390 2.480 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.315  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.520 16.440 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 29.120 5.600 ;
        RECT  28.420 4.610 28.820 5.600 ;
        RECT  27.120 4.620 27.520 5.600 ;
        RECT  25.700 4.610 26.100 5.600 ;
        RECT  24.400 4.620 24.800 5.600 ;
        RECT  23.090 4.620 23.490 5.600 ;
        RECT  19.740 4.710 20.140 5.600 ;
        RECT  17.750 4.340 17.990 5.600 ;
        RECT  15.850 4.340 16.090 5.600 ;
        RECT  13.690 4.710 14.090 5.600 ;
        RECT  9.370 4.710 9.780 5.600 ;
        RECT  8.190 4.710 8.590 5.600 ;
        RECT  2.940 3.950 3.180 5.600 ;
        RECT  0.730 4.710 1.130 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 29.120 0.740 ;
        RECT  28.330 0.000 28.730 0.890 ;
        RECT  26.970 0.000 27.370 0.890 ;
        RECT  25.610 0.000 26.010 0.890 ;
        RECT  24.250 0.000 24.650 0.890 ;
        RECT  22.890 0.000 23.290 0.890 ;
        RECT  18.410 0.000 18.810 0.890 ;
        RECT  17.290 0.000 17.690 0.820 ;
        RECT  16.350 0.000 16.590 1.260 ;
        RECT  9.460 0.000 9.860 0.890 ;
        RECT  8.600 0.000 9.000 0.890 ;
        RECT  3.120 0.000 3.520 0.940 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.180 2.090 ;
        RECT  0.940 2.470 1.510 2.870 ;
        RECT  0.940 1.850 1.180 3.650 ;
        RECT  0.150 3.410 1.180 3.650 ;
        RECT  1.590 1.770 1.990 2.170 ;
        RECT  1.750 2.600 2.620 2.840 ;
        RECT  1.750 1.770 1.990 3.500 ;
        RECT  1.590 3.100 1.990 3.500 ;
        RECT  2.290 3.330 3.670 3.570 ;
        RECT  3.430 3.330 3.670 3.940 ;
        RECT  3.430 3.700 5.660 3.940 ;
        RECT  3.920 0.980 5.790 1.220 ;
        RECT  6.240 0.980 8.040 1.220 ;
        RECT  4.620 1.470 5.850 1.710 ;
        RECT  5.610 1.470 5.850 1.970 ;
        RECT  6.240 0.980 6.480 1.970 ;
        RECT  5.610 1.730 6.480 1.970 ;
        RECT  7.980 1.750 8.840 1.990 ;
        RECT  7.980 1.750 8.220 3.390 ;
        RECT  7.390 3.060 8.220 3.390 ;
        RECT  7.390 3.060 7.800 3.990 ;
        RECT  7.060 3.750 7.800 3.990 ;
        RECT  10.620 1.460 11.560 1.700 ;
        RECT  10.620 1.460 11.030 1.860 ;
        RECT  10.620 1.460 10.950 2.530 ;
        RECT  10.230 2.290 10.950 2.530 ;
        RECT  10.230 2.290 10.470 3.990 ;
        RECT  10.230 3.750 11.080 3.990 ;
        RECT  1.890 1.150 2.860 1.390 ;
        RECT  2.620 1.150 2.860 1.700 ;
        RECT  2.620 1.460 4.300 1.700 ;
        RECT  6.740 1.540 7.300 1.780 ;
        RECT  11.820 1.770 12.060 2.440 ;
        RECT  11.210 2.200 12.060 2.440 ;
        RECT  4.060 1.460 4.300 3.460 ;
        RECT  6.740 1.540 6.980 3.470 ;
        RECT  11.210 2.200 11.620 3.450 ;
        RECT  4.060 3.040 7.100 3.460 ;
        RECT  6.440 3.040 7.100 3.470 ;
        RECT  6.440 3.040 6.680 4.470 ;
        RECT  11.380 2.200 11.620 4.470 ;
        RECT  6.440 4.230 11.620 4.470 ;
        RECT  13.150 1.550 13.830 1.790 ;
        RECT  13.150 1.550 13.390 2.380 ;
        RECT  12.780 2.140 13.390 2.380 ;
        RECT  12.780 2.140 13.020 3.390 ;
        RECT  12.780 3.150 13.850 3.390 ;
        RECT  13.610 3.300 14.690 3.540 ;
        RECT  12.300 1.580 12.910 1.820 ;
        RECT  12.300 1.580 12.540 3.090 ;
        RECT  11.860 2.850 12.540 3.090 ;
        RECT  11.860 2.850 12.100 4.390 ;
        RECT  11.860 4.150 15.610 4.390 ;
        RECT  17.580 2.170 19.790 2.410 ;
        RECT  17.580 1.770 17.820 3.370 ;
        RECT  17.080 3.130 18.890 3.370 ;
        RECT  10.130 0.980 16.030 1.220 ;
        RECT  19.200 0.980 21.080 1.220 ;
        RECT  16.940 1.130 19.440 1.370 ;
        RECT  15.790 0.980 16.030 1.740 ;
        RECT  16.940 1.130 17.180 1.740 ;
        RECT  15.790 1.500 17.180 1.740 ;
        RECT  10.130 0.980 10.370 2.050 ;
        RECT  9.150 1.810 10.370 2.050 ;
        RECT  9.740 1.810 9.980 3.990 ;
        RECT  8.700 3.750 9.980 3.990 ;
        RECT  18.060 1.620 20.270 1.860 ;
        RECT  20.030 1.620 20.270 3.510 ;
        RECT  19.550 3.130 20.270 3.370 ;
        RECT  20.030 3.270 21.310 3.510 ;
        RECT  21.800 1.850 22.450 2.090 ;
        RECT  15.070 1.770 15.510 2.180 ;
        RECT  13.630 2.040 15.310 2.280 ;
        RECT  13.630 2.040 13.870 2.860 ;
        RECT  13.260 2.620 13.870 2.860 ;
        RECT  22.210 1.850 22.450 3.580 ;
        RECT  14.990 2.040 15.310 3.660 ;
        RECT  22.210 3.170 22.800 3.580 ;
        RECT  14.990 3.260 16.780 3.660 ;
        RECT  16.450 3.610 18.700 3.850 ;
        RECT  18.460 3.610 18.700 4.470 ;
        RECT  22.470 3.170 22.800 4.470 ;
        RECT  18.460 4.230 22.800 4.470 ;
        RECT  21.270 1.370 22.930 1.610 ;
        RECT  20.910 1.550 21.510 1.960 ;
        RECT  22.690 1.370 22.930 2.860 ;
        RECT  20.910 1.550 21.230 2.800 ;
        RECT  20.910 2.560 21.970 2.800 ;
        RECT  22.690 2.460 23.320 2.860 ;
        RECT  19.020 3.610 19.790 3.850 ;
        RECT  21.730 2.560 21.970 3.990 ;
        RECT  19.550 3.750 21.970 3.990 ;
    END
END skbrb4

MACRO skbrb2
    CLASS CORE ;
    FOREIGN skbrb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.320 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.110 2.520 14.660 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.243  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 2.580 9.350 3.160 ;
        END
    END CP
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.369  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 5.070 2.480 ;
        END
    END J
    PIN KZ
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.020 7.740 2.600 ;
        END
    END KZ
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.283  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  24.960 2.580 25.420 4.180 ;
        RECT  25.020 1.770 25.420 4.180 ;
        RECT  24.700 2.580 25.420 3.020 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.285  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  23.660 1.770 24.060 4.150 ;
        RECT  23.570 2.530 24.060 3.020 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.700 3.130 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.390 2.480 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.315  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.520 16.440 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 26.320 5.600 ;
        RECT  25.700 4.610 26.100 5.600 ;
        RECT  24.400 4.620 24.800 5.600 ;
        RECT  23.090 4.620 23.490 5.600 ;
        RECT  19.740 4.710 20.140 5.600 ;
        RECT  17.750 4.340 17.990 5.600 ;
        RECT  15.850 4.340 16.090 5.600 ;
        RECT  13.690 4.710 14.090 5.600 ;
        RECT  9.370 4.710 9.780 5.600 ;
        RECT  8.190 4.710 8.590 5.600 ;
        RECT  2.940 3.950 3.180 5.600 ;
        RECT  0.730 4.710 1.130 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 26.320 0.740 ;
        RECT  25.610 0.000 26.010 0.890 ;
        RECT  24.250 0.000 24.650 0.890 ;
        RECT  22.890 0.000 23.290 0.890 ;
        RECT  18.410 0.000 18.810 0.890 ;
        RECT  17.330 0.000 17.730 0.820 ;
        RECT  16.350 0.000 16.590 1.260 ;
        RECT  9.460 0.000 9.860 0.890 ;
        RECT  8.600 0.000 9.000 0.890 ;
        RECT  3.120 0.000 3.520 0.940 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.180 2.090 ;
        RECT  0.940 2.470 1.510 2.870 ;
        RECT  0.940 1.850 1.180 3.650 ;
        RECT  0.150 3.410 1.180 3.650 ;
        RECT  1.590 1.770 1.990 2.170 ;
        RECT  1.750 2.600 2.620 2.840 ;
        RECT  1.750 1.770 1.990 3.500 ;
        RECT  1.590 3.100 1.990 3.500 ;
        RECT  2.290 3.330 3.660 3.570 ;
        RECT  3.420 3.330 3.660 3.940 ;
        RECT  3.420 3.700 5.660 3.940 ;
        RECT  3.920 0.980 5.790 1.220 ;
        RECT  6.240 0.980 8.040 1.220 ;
        RECT  4.620 1.470 5.850 1.710 ;
        RECT  5.610 1.470 5.850 1.970 ;
        RECT  6.240 0.980 6.480 1.970 ;
        RECT  5.610 1.730 6.480 1.970 ;
        RECT  7.980 1.750 8.840 1.990 ;
        RECT  7.980 1.750 8.220 3.390 ;
        RECT  7.390 3.060 8.220 3.390 ;
        RECT  7.390 3.060 7.720 3.990 ;
        RECT  7.060 3.750 7.720 3.990 ;
        RECT  10.620 1.460 11.560 1.700 ;
        RECT  10.620 1.460 11.030 1.860 ;
        RECT  10.620 1.460 10.950 2.530 ;
        RECT  10.230 2.290 10.950 2.530 ;
        RECT  10.230 2.290 10.470 3.990 ;
        RECT  10.230 3.750 11.080 3.990 ;
        RECT  1.890 1.150 2.860 1.390 ;
        RECT  2.620 1.150 2.860 1.700 ;
        RECT  2.620 1.460 4.300 1.700 ;
        RECT  6.740 1.540 7.300 1.780 ;
        RECT  11.820 1.770 12.060 2.520 ;
        RECT  11.210 2.280 12.060 2.520 ;
        RECT  4.060 1.460 4.300 3.460 ;
        RECT  6.740 1.540 6.980 3.470 ;
        RECT  11.210 2.280 11.620 3.450 ;
        RECT  4.060 3.040 6.980 3.460 ;
        RECT  6.500 3.070 7.100 3.470 ;
        RECT  6.500 3.040 6.740 4.470 ;
        RECT  11.380 2.280 11.620 4.470 ;
        RECT  6.500 4.230 11.620 4.470 ;
        RECT  13.150 1.460 13.760 1.700 ;
        RECT  13.150 1.460 13.390 2.380 ;
        RECT  12.780 2.140 13.390 2.380 ;
        RECT  12.780 2.140 13.020 3.390 ;
        RECT  12.780 3.150 13.850 3.390 ;
        RECT  13.610 3.300 14.690 3.540 ;
        RECT  12.300 1.580 12.910 1.820 ;
        RECT  12.300 1.580 12.540 3.090 ;
        RECT  11.860 2.850 12.540 3.090 ;
        RECT  11.860 2.850 12.100 4.390 ;
        RECT  11.860 4.150 15.610 4.390 ;
        RECT  17.580 2.170 19.790 2.410 ;
        RECT  17.580 1.770 17.820 3.370 ;
        RECT  17.080 3.130 18.890 3.370 ;
        RECT  10.130 0.980 16.030 1.220 ;
        RECT  19.170 0.980 21.080 1.220 ;
        RECT  16.940 1.130 19.410 1.370 ;
        RECT  15.790 0.980 16.030 1.740 ;
        RECT  16.940 1.130 17.180 1.740 ;
        RECT  15.790 1.500 17.180 1.740 ;
        RECT  10.130 0.980 10.370 2.050 ;
        RECT  9.150 1.810 10.370 2.050 ;
        RECT  9.740 1.810 9.980 3.990 ;
        RECT  8.700 3.750 9.980 3.990 ;
        RECT  18.060 1.620 20.270 1.860 ;
        RECT  20.030 1.620 20.270 3.510 ;
        RECT  19.550 3.130 20.270 3.370 ;
        RECT  20.030 3.270 21.310 3.510 ;
        RECT  21.800 1.850 22.450 2.090 ;
        RECT  15.070 1.770 15.510 2.180 ;
        RECT  13.630 2.030 15.390 2.270 ;
        RECT  13.630 2.030 13.870 2.860 ;
        RECT  13.260 2.620 13.870 2.860 ;
        RECT  22.210 1.850 22.450 3.580 ;
        RECT  14.980 2.030 15.390 3.660 ;
        RECT  22.210 3.170 22.800 3.580 ;
        RECT  14.980 3.260 16.780 3.660 ;
        RECT  16.450 3.610 18.670 3.850 ;
        RECT  18.430 3.610 18.670 4.470 ;
        RECT  22.470 3.170 22.800 4.470 ;
        RECT  18.430 4.230 22.800 4.470 ;
        RECT  21.270 1.370 22.930 1.610 ;
        RECT  20.910 1.550 21.510 1.960 ;
        RECT  22.690 1.370 22.930 2.860 ;
        RECT  20.910 1.550 21.230 2.800 ;
        RECT  20.910 2.560 21.970 2.800 ;
        RECT  22.690 2.460 23.320 2.860 ;
        RECT  19.020 3.610 19.790 3.850 ;
        RECT  21.730 2.560 21.970 3.990 ;
        RECT  19.550 3.750 21.970 3.990 ;
    END
END skbrb2

MACRO skbrb1
    CLASS CORE ;
    FOREIGN skbrb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.060 2.520 14.690 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.243  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 2.580 9.350 3.160 ;
        END
    END CP
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.369  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 5.070 2.480 ;
        END
    END J
    PIN KZ
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.020 7.740 2.600 ;
        END
    END KZ
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  24.670 1.770 25.080 3.490 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.313  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  23.090 2.530 24.020 3.020 ;
        RECT  23.090 1.770 23.490 4.000 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.700 3.130 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.390 2.480 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.315  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.520 16.440 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 25.200 5.600 ;
        RECT  23.760 4.710 24.160 5.600 ;
        RECT  19.740 4.710 20.140 5.600 ;
        RECT  17.750 4.340 17.990 5.600 ;
        RECT  15.850 4.340 16.090 5.600 ;
        RECT  13.690 4.710 14.090 5.600 ;
        RECT  9.370 4.710 9.780 5.600 ;
        RECT  8.190 4.710 8.590 5.600 ;
        RECT  2.940 3.950 3.180 5.600 ;
        RECT  0.730 4.710 1.140 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 25.200 0.740 ;
        RECT  23.820 0.000 24.220 0.890 ;
        RECT  18.410 0.000 18.810 0.890 ;
        RECT  17.370 0.000 17.770 0.820 ;
        RECT  16.350 0.000 16.590 1.260 ;
        RECT  9.460 0.000 9.860 0.890 ;
        RECT  8.600 0.000 9.000 0.890 ;
        RECT  3.120 0.000 3.520 0.940 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.180 2.090 ;
        RECT  0.940 2.520 1.510 2.920 ;
        RECT  0.940 1.850 1.180 3.650 ;
        RECT  0.150 3.410 1.180 3.650 ;
        RECT  1.590 1.770 2.000 2.170 ;
        RECT  1.760 2.600 2.620 2.840 ;
        RECT  1.760 1.770 2.000 3.550 ;
        RECT  1.590 3.150 2.000 3.550 ;
        RECT  2.290 3.330 3.820 3.570 ;
        RECT  3.580 3.330 3.820 3.940 ;
        RECT  3.580 3.700 5.660 3.940 ;
        RECT  3.920 0.980 5.790 1.220 ;
        RECT  6.240 0.980 8.040 1.220 ;
        RECT  4.620 1.470 5.850 1.710 ;
        RECT  5.610 1.470 5.850 1.970 ;
        RECT  6.240 0.980 6.480 1.970 ;
        RECT  5.610 1.730 6.480 1.970 ;
        RECT  7.980 1.750 8.840 1.990 ;
        RECT  7.980 1.750 8.220 3.150 ;
        RECT  7.480 2.910 8.220 3.150 ;
        RECT  7.480 2.910 7.720 3.990 ;
        RECT  7.060 3.750 7.720 3.990 ;
        RECT  10.630 1.460 11.560 1.700 ;
        RECT  10.630 1.460 11.030 1.850 ;
        RECT  10.630 1.460 10.950 2.530 ;
        RECT  10.230 2.290 10.950 2.530 ;
        RECT  10.230 2.290 10.470 3.990 ;
        RECT  10.230 3.750 11.080 3.990 ;
        RECT  1.890 1.150 2.860 1.390 ;
        RECT  2.620 1.150 2.860 1.700 ;
        RECT  2.620 1.460 4.300 1.700 ;
        RECT  6.740 1.540 7.300 1.780 ;
        RECT  11.800 1.700 12.040 2.370 ;
        RECT  11.210 2.130 12.040 2.370 ;
        RECT  4.060 1.460 4.300 3.450 ;
        RECT  6.740 1.540 6.980 3.480 ;
        RECT  4.060 3.050 7.100 3.450 ;
        RECT  11.210 2.130 11.450 3.450 ;
        RECT  6.580 3.050 7.100 3.480 ;
        RECT  6.580 3.050 6.820 4.470 ;
        RECT  11.380 3.050 11.620 4.470 ;
        RECT  6.580 4.230 11.620 4.470 ;
        RECT  13.100 1.460 13.760 1.700 ;
        RECT  13.100 1.460 13.340 2.380 ;
        RECT  12.780 2.140 13.340 2.380 ;
        RECT  12.780 2.140 13.020 3.390 ;
        RECT  12.780 3.150 13.850 3.390 ;
        RECT  13.610 3.300 14.690 3.540 ;
        RECT  12.280 1.660 12.860 1.900 ;
        RECT  12.280 1.660 12.520 3.090 ;
        RECT  11.860 2.850 12.520 3.090 ;
        RECT  11.860 2.850 12.100 4.530 ;
        RECT  12.370 4.150 15.610 4.390 ;
        RECT  11.860 4.290 12.600 4.530 ;
        RECT  17.580 2.170 19.790 2.410 ;
        RECT  17.580 1.770 17.820 3.370 ;
        RECT  17.080 3.130 18.890 3.370 ;
        RECT  10.100 0.980 16.030 1.220 ;
        RECT  19.190 0.980 21.080 1.220 ;
        RECT  16.940 1.130 19.430 1.370 ;
        RECT  15.790 0.980 16.030 1.740 ;
        RECT  10.100 0.980 10.340 1.510 ;
        RECT  16.940 1.130 17.180 1.740 ;
        RECT  15.790 1.500 17.180 1.740 ;
        RECT  9.970 1.270 10.230 2.050 ;
        RECT  9.150 1.810 10.230 2.050 ;
        RECT  9.740 1.810 9.980 3.990 ;
        RECT  8.700 3.750 9.980 3.990 ;
        RECT  18.060 1.620 20.270 1.860 ;
        RECT  20.030 1.620 20.270 3.510 ;
        RECT  19.550 3.130 20.270 3.370 ;
        RECT  20.030 3.270 21.310 3.510 ;
        RECT  21.800 1.640 22.710 1.880 ;
        RECT  15.070 1.770 15.510 2.180 ;
        RECT  13.580 1.940 15.510 2.180 ;
        RECT  13.580 1.940 13.820 2.860 ;
        RECT  13.260 2.620 13.820 2.860 ;
        RECT  15.020 1.940 15.420 3.590 ;
        RECT  15.020 3.270 16.780 3.590 ;
        RECT  16.370 3.270 16.780 3.850 ;
        RECT  16.370 3.610 18.550 3.850 ;
        RECT  18.310 3.610 18.550 4.470 ;
        RECT  22.470 1.640 22.710 4.470 ;
        RECT  18.310 4.230 22.710 4.470 ;
        RECT  21.320 1.050 23.630 1.290 ;
        RECT  21.320 1.050 21.560 1.950 ;
        RECT  20.910 1.560 21.560 1.950 ;
        RECT  20.910 1.560 21.230 2.800 ;
        RECT  20.910 2.560 21.970 2.800 ;
        RECT  19.020 3.610 19.680 3.850 ;
        RECT  21.730 2.560 21.970 3.990 ;
        RECT  19.460 3.750 21.970 3.990 ;
    END
END skbrb1

MACRO seprq4
    CLASS CORE ;
    FOREIGN seprq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 23.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.516  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 2.580 9.520 3.020 ;
        RECT  9.280 2.180 9.520 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.230 1.680 4.980 1.920 ;
        RECT  4.540 1.460 4.980 1.920 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.899  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.570 2.950 5.780 3.190 ;
        RECT  5.540 2.630 5.780 3.190 ;
        RECT  2.860 2.870 4.760 3.110 ;
        RECT  2.860 2.580 3.300 3.110 ;
        RECT  2.860 2.180 3.220 3.110 ;
        RECT  2.820 2.180 3.220 2.540 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.125  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.470 3.150 19.590 3.390 ;
        RECT  18.020 1.850 19.340 2.090 ;
        RECT  17.470 2.370 18.260 2.610 ;
        RECT  17.980 2.020 18.420 2.460 ;
        RECT  17.470 1.770 17.710 3.390 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.529  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.230 2.510 0.630 2.940 ;
        RECT  0.120 2.580 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.369  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.020 7.630 2.460 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.600 2.520 14.000 2.900 ;
        RECT  13.500 2.580 13.940 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 23.520 5.600 ;
        RECT  19.740 4.610 20.140 5.600 ;
        RECT  18.450 4.610 18.850 5.600 ;
        RECT  17.130 4.620 17.530 5.600 ;
        RECT  15.750 3.870 15.990 5.600 ;
        RECT  14.410 4.710 14.810 5.600 ;
        RECT  13.010 4.710 13.410 5.600 ;
        RECT  11.170 4.780 11.570 5.600 ;
        RECT  9.620 4.610 10.020 5.600 ;
        RECT  6.490 3.980 6.730 5.600 ;
        RECT  2.950 4.140 3.190 5.600 ;
        RECT  0.900 4.380 1.300 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 23.520 0.740 ;
        RECT  19.710 0.000 20.110 1.260 ;
        RECT  18.170 0.000 18.570 1.260 ;
        RECT  15.310 0.000 15.550 1.650 ;
        RECT  13.340 0.000 13.580 1.640 ;
        RECT  9.470 0.000 9.870 0.890 ;
        RECT  7.050 0.000 7.290 1.220 ;
        RECT  2.790 0.000 3.200 0.890 ;
        RECT  0.920 0.000 1.320 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.140 1.450 1.230 1.690 ;
        RECT  0.990 1.450 1.230 4.030 ;
        RECT  0.140 3.790 1.230 4.030 ;
        RECT  1.590 1.510 1.830 2.480 ;
        RECT  1.780 2.240 2.020 3.200 ;
        RECT  1.550 2.960 1.790 3.510 ;
        RECT  2.210 1.480 2.530 1.810 ;
        RECT  2.210 1.570 3.870 1.810 ;
        RECT  3.630 1.570 3.870 2.590 ;
        RECT  2.290 1.480 2.530 3.260 ;
        RECT  2.380 2.990 2.620 3.710 ;
        RECT  5.480 1.740 5.720 2.390 ;
        RECT  5.060 2.150 6.310 2.390 ;
        RECT  5.480 2.140 6.310 2.390 ;
        RECT  4.250 2.360 5.300 2.600 ;
        RECT  6.070 2.140 6.310 3.000 ;
        RECT  8.020 2.430 8.260 3.000 ;
        RECT  6.070 2.760 8.260 3.000 ;
        RECT  8.980 1.680 10.010 1.920 ;
        RECT  9.770 2.290 10.330 2.530 ;
        RECT  9.770 1.680 10.010 3.890 ;
        RECT  9.040 3.650 10.010 3.890 ;
        RECT  10.340 1.650 10.870 2.050 ;
        RECT  10.630 2.280 11.010 2.680 ;
        RECT  10.630 1.650 10.870 3.020 ;
        RECT  10.440 2.780 10.680 3.550 ;
        RECT  4.500 0.980 6.560 1.220 ;
        RECT  10.340 1.010 11.360 1.250 ;
        RECT  7.660 1.170 10.580 1.410 ;
        RECT  6.320 0.980 6.560 1.740 ;
        RECT  7.660 1.170 7.900 1.740 ;
        RECT  6.320 1.500 7.900 1.740 ;
        RECT  11.120 1.010 11.360 1.880 ;
        RECT  11.300 1.640 11.540 3.150 ;
        RECT  6.070 3.240 8.740 3.480 ;
        RECT  8.500 1.170 8.740 3.480 ;
        RECT  11.140 2.910 11.380 3.480 ;
        RECT  4.630 3.470 6.320 3.740 ;
        RECT  4.630 3.470 4.870 4.570 ;
        RECT  12.470 1.250 12.920 1.650 ;
        RECT  12.470 1.250 12.710 3.480 ;
        RECT  11.780 1.500 12.230 1.900 ;
        RECT  11.990 1.500 12.230 3.990 ;
        RECT  11.990 3.750 14.660 3.990 ;
        RECT  14.420 2.390 14.660 3.990 ;
        RECT  11.640 3.810 12.170 4.050 ;
        RECT  19.960 2.250 20.800 2.490 ;
        RECT  20.560 1.620 20.800 2.490 ;
        RECT  18.660 2.430 20.210 2.670 ;
        RECT  19.970 2.250 20.210 3.380 ;
        RECT  19.970 3.140 20.940 3.380 ;
        RECT  15.920 1.010 17.230 1.250 ;
        RECT  14.610 1.570 14.850 2.140 ;
        RECT  15.920 1.010 16.160 2.140 ;
        RECT  13.000 1.900 16.160 2.140 ;
        RECT  21.260 0.980 21.500 2.760 ;
        RECT  21.260 2.520 21.850 2.760 ;
        RECT  13.000 1.900 13.240 3.500 ;
        RECT  13.000 3.260 14.180 3.500 ;
        RECT  16.990 1.010 17.230 3.870 ;
        RECT  21.260 3.410 21.850 3.650 ;
        RECT  21.610 2.520 21.850 3.650 ;
        RECT  16.990 3.630 21.500 3.870 ;
        RECT  21.920 0.980 22.420 1.380 ;
        RECT  22.180 0.980 22.420 3.320 ;
        RECT  22.270 3.070 22.510 4.130 ;
        RECT  21.910 3.890 22.510 4.130 ;
        RECT  22.660 0.980 23.010 1.380 ;
        RECT  16.510 1.650 16.750 2.820 ;
        RECT  15.180 2.580 16.750 2.820 ;
        RECT  16.500 2.580 16.740 4.350 ;
        RECT  12.390 4.230 15.420 4.470 ;
        RECT  16.500 4.110 21.500 4.350 ;
        RECT  9.040 4.130 10.680 4.370 ;
        RECT  21.260 4.110 21.500 4.620 ;
        RECT  15.180 2.580 15.420 4.470 ;
        RECT  10.440 4.300 12.690 4.540 ;
        RECT  9.040 4.130 9.280 4.620 ;
        RECT  8.080 4.380 9.280 4.620 ;
        RECT  22.770 0.980 23.010 4.620 ;
        RECT  21.260 4.380 23.010 4.620 ;
    END
END seprq4

MACRO seprq2
    CLASS CORE ;
    FOREIGN seprq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 28.560 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.580 16.630 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.940 2.250 13.380 3.020 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.397  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.700 2.580 7.310 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.159  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  26.940 3.110 27.830 3.580 ;
        RECT  27.510 1.240 27.830 3.580 ;
        RECT  27.430 1.240 27.830 1.640 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.020 0.980 2.900 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.280 1.640 3.020 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.241  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  25.260 2.190 25.720 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 28.560 5.600 ;
        RECT  28.070 4.190 28.310 5.600 ;
        RECT  26.770 4.190 27.010 5.600 ;
        RECT  25.860 4.390 26.260 5.600 ;
        RECT  24.380 4.390 24.780 5.600 ;
        RECT  21.610 4.710 22.010 5.600 ;
        RECT  20.420 4.710 20.820 5.600 ;
        RECT  16.580 4.640 16.980 5.600 ;
        RECT  14.770 4.330 15.010 5.600 ;
        RECT  13.390 4.710 13.790 5.600 ;
        RECT  9.670 4.480 10.070 5.600 ;
        RECT  8.200 3.770 8.440 5.600 ;
        RECT  6.900 3.770 7.140 5.600 ;
        RECT  6.000 3.850 6.240 5.600 ;
        RECT  3.930 4.090 4.170 5.600 ;
        RECT  1.660 4.460 2.060 5.600 ;
        RECT  0.970 3.290 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 28.560 0.740 ;
        RECT  28.010 0.000 28.410 0.980 ;
        RECT  26.660 0.000 27.060 0.980 ;
        RECT  25.260 0.000 25.500 1.380 ;
        RECT  20.550 0.000 20.790 1.830 ;
        RECT  16.750 0.000 17.150 0.890 ;
        RECT  15.420 0.000 15.820 0.890 ;
        RECT  13.210 0.000 13.610 0.890 ;
        RECT  10.240 0.000 10.640 0.890 ;
        RECT  8.130 0.000 8.530 0.890 ;
        RECT  6.180 0.000 6.600 0.890 ;
        RECT  4.190 0.000 4.430 1.470 ;
        RECT  1.660 0.000 2.060 1.140 ;
        RECT  0.760 0.000 1.180 1.180 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 1.520 0.470 1.920 ;
        RECT  0.220 1.520 0.460 4.620 ;
        RECT  0.220 3.290 0.470 4.620 ;
        RECT  1.570 1.530 2.120 1.930 ;
        RECT  1.880 2.270 2.990 2.510 ;
        RECT  1.880 1.530 2.120 3.650 ;
        RECT  1.630 3.260 2.120 3.650 ;
        RECT  2.430 0.980 2.990 1.380 ;
        RECT  2.670 0.980 2.990 1.910 ;
        RECT  2.670 1.630 3.470 1.910 ;
        RECT  3.230 1.630 3.470 2.990 ;
        RECT  2.480 2.750 3.470 2.990 ;
        RECT  2.480 2.750 2.720 4.620 ;
        RECT  2.430 4.220 2.830 4.620 ;
        RECT  3.230 1.150 3.950 1.390 ;
        RECT  3.710 2.800 4.450 3.040 ;
        RECT  3.710 1.150 3.950 3.610 ;
        RECT  2.960 3.370 3.950 3.610 ;
        RECT  2.960 3.370 3.360 3.770 ;
        RECT  4.570 1.830 4.930 2.230 ;
        RECT  4.690 1.830 4.930 3.750 ;
        RECT  4.430 3.350 4.930 3.750 ;
        RECT  6.000 1.610 6.580 1.850 ;
        RECT  6.000 1.610 6.240 3.510 ;
        RECT  9.440 1.610 9.680 2.500 ;
        RECT  9.160 2.260 10.350 2.500 ;
        RECT  9.160 2.260 9.400 3.740 ;
        RECT  10.240 1.690 10.890 1.930 ;
        RECT  10.650 2.510 11.050 2.910 ;
        RECT  10.650 1.690 10.890 3.740 ;
        RECT  10.440 3.340 10.890 3.740 ;
        RECT  12.460 1.610 13.020 2.010 ;
        RECT  12.460 1.610 12.700 3.510 ;
        RECT  12.460 3.270 13.020 3.510 ;
        RECT  6.900 1.620 7.860 1.860 ;
        RECT  7.620 1.620 7.860 3.510 ;
        RECT  7.540 3.110 7.940 3.510 ;
        RECT  7.540 3.270 8.920 3.510 ;
        RECT  8.680 3.270 8.920 4.240 ;
        RECT  8.680 4.000 10.600 4.240 ;
        RECT  10.360 4.000 10.600 4.530 ;
        RECT  12.900 4.230 14.140 4.470 ;
        RECT  10.360 4.290 13.140 4.530 ;
        RECT  14.070 2.140 14.670 2.540 ;
        RECT  14.070 1.610 14.310 3.510 ;
        RECT  11.140 1.610 11.540 2.010 ;
        RECT  11.300 1.610 11.540 4.050 ;
        RECT  11.140 3.250 11.540 4.050 ;
        RECT  14.750 3.590 15.150 3.990 ;
        RECT  12.400 3.750 15.150 3.990 ;
        RECT  14.910 1.610 15.150 3.990 ;
        RECT  11.140 3.810 12.700 4.050 ;
        RECT  16.120 1.860 17.110 2.100 ;
        RECT  16.870 2.360 17.500 2.600 ;
        RECT  16.870 1.860 17.110 3.530 ;
        RECT  16.050 3.290 17.110 3.530 ;
        RECT  5.390 1.130 18.500 1.370 ;
        RECT  18.220 1.130 18.500 3.510 ;
        RECT  11.960 1.130 12.200 3.570 ;
        RECT  5.390 1.130 5.630 3.650 ;
        RECT  5.170 3.250 5.630 3.650 ;
        RECT  17.480 1.720 17.980 2.120 ;
        RECT  17.350 3.290 17.980 3.530 ;
        RECT  17.740 1.720 17.980 4.060 ;
        RECT  17.740 3.820 18.760 4.060 ;
        RECT  19.660 1.450 20.060 1.850 ;
        RECT  19.720 1.450 19.960 3.510 ;
        RECT  19.600 3.110 20.020 3.510 ;
        RECT  18.880 3.110 19.280 3.510 ;
        RECT  19.000 1.450 19.240 3.990 ;
        RECT  21.590 2.580 21.830 3.990 ;
        RECT  19.000 3.750 21.830 3.990 ;
        RECT  20.200 2.100 22.630 2.340 ;
        RECT  21.080 2.100 21.320 3.510 ;
        RECT  22.390 1.640 22.630 3.720 ;
        RECT  15.390 3.840 15.790 4.370 ;
        RECT  23.870 3.910 25.440 4.150 ;
        RECT  18.930 4.230 24.110 4.470 ;
        RECT  15.390 4.130 17.460 4.370 ;
        RECT  23.870 1.640 24.110 4.470 ;
        RECT  17.220 4.300 19.100 4.540 ;
        RECT  25.200 3.910 25.440 4.620 ;
        RECT  23.130 1.160 24.590 1.400 ;
        RECT  24.350 1.160 24.590 1.940 ;
        RECT  24.350 1.700 26.200 1.940 ;
        RECT  25.960 1.840 26.540 2.090 ;
        RECT  23.130 1.160 23.370 3.720 ;
        RECT  25.880 1.220 27.020 1.460 ;
        RECT  26.780 1.220 27.020 2.570 ;
        RECT  26.780 2.170 27.270 2.570 ;
        RECT  26.050 2.330 27.270 2.570 ;
        RECT  24.870 3.270 26.290 3.510 ;
        RECT  26.050 2.330 26.290 3.670 ;
        RECT  25.890 3.270 26.290 3.670 ;
    END
END seprq2

MACRO seprq1
    CLASS CORE ;
    FOREIGN seprq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 28.000 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.580 16.630 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.940 2.250 13.380 3.020 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.397  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.700 2.580 7.310 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.264  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  26.940 3.110 27.830 3.580 ;
        RECT  27.510 1.240 27.830 3.580 ;
        RECT  27.430 1.240 27.830 1.640 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.020 0.980 2.900 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.280 1.640 3.020 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.241  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  25.260 2.190 25.720 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 28.000 5.600 ;
        RECT  26.770 4.190 27.010 5.600 ;
        RECT  25.860 4.390 26.260 5.600 ;
        RECT  24.380 4.390 24.780 5.600 ;
        RECT  21.610 4.710 22.010 5.600 ;
        RECT  20.420 4.710 20.820 5.600 ;
        RECT  16.580 4.640 16.980 5.600 ;
        RECT  14.770 4.330 15.010 5.600 ;
        RECT  13.390 4.710 13.790 5.600 ;
        RECT  9.670 4.480 10.070 5.600 ;
        RECT  8.200 3.770 8.440 5.600 ;
        RECT  6.900 3.770 7.140 5.600 ;
        RECT  6.000 3.850 6.240 5.600 ;
        RECT  3.930 4.090 4.170 5.600 ;
        RECT  1.660 4.460 2.060 5.600 ;
        RECT  0.970 3.290 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 28.000 0.740 ;
        RECT  26.660 0.000 27.060 0.980 ;
        RECT  25.260 0.000 25.500 1.380 ;
        RECT  20.550 0.000 20.790 1.830 ;
        RECT  16.750 0.000 17.150 0.890 ;
        RECT  15.420 0.000 15.820 0.890 ;
        RECT  13.210 0.000 13.610 0.890 ;
        RECT  10.240 0.000 10.640 0.890 ;
        RECT  8.130 0.000 8.530 0.890 ;
        RECT  6.180 0.000 6.600 0.890 ;
        RECT  4.190 0.000 4.430 1.470 ;
        RECT  1.660 0.000 2.060 1.140 ;
        RECT  0.760 0.000 1.180 1.180 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 1.520 0.470 1.920 ;
        RECT  0.220 1.520 0.460 4.620 ;
        RECT  0.220 3.290 0.470 4.620 ;
        RECT  1.570 1.530 2.120 1.930 ;
        RECT  1.880 2.270 2.990 2.510 ;
        RECT  1.880 1.530 2.120 3.650 ;
        RECT  1.630 3.260 2.120 3.650 ;
        RECT  2.430 0.980 2.990 1.380 ;
        RECT  2.670 0.980 2.990 1.910 ;
        RECT  2.670 1.630 3.470 1.910 ;
        RECT  3.230 1.630 3.470 2.990 ;
        RECT  2.480 2.750 3.470 2.990 ;
        RECT  2.480 2.750 2.720 4.620 ;
        RECT  2.430 4.220 2.830 4.620 ;
        RECT  3.230 1.150 3.950 1.390 ;
        RECT  3.710 2.800 4.450 3.040 ;
        RECT  3.710 1.150 3.950 3.610 ;
        RECT  2.960 3.370 3.950 3.610 ;
        RECT  2.960 3.370 3.360 3.770 ;
        RECT  4.570 1.830 4.930 2.230 ;
        RECT  4.690 1.830 4.930 3.750 ;
        RECT  4.430 3.350 4.930 3.750 ;
        RECT  6.000 1.610 6.580 1.850 ;
        RECT  6.000 1.610 6.240 3.510 ;
        RECT  9.440 1.610 9.680 2.500 ;
        RECT  9.160 2.260 10.350 2.500 ;
        RECT  9.160 2.260 9.400 3.740 ;
        RECT  10.240 1.690 10.890 1.930 ;
        RECT  10.650 2.510 11.050 2.910 ;
        RECT  10.650 1.690 10.890 3.740 ;
        RECT  10.440 3.340 10.890 3.740 ;
        RECT  12.460 1.610 13.020 2.010 ;
        RECT  12.460 1.610 12.700 3.510 ;
        RECT  12.460 3.270 13.020 3.510 ;
        RECT  6.900 1.620 7.860 1.860 ;
        RECT  7.620 1.620 7.860 3.510 ;
        RECT  7.540 3.110 7.940 3.510 ;
        RECT  7.540 3.270 8.920 3.510 ;
        RECT  8.680 3.270 8.920 4.240 ;
        RECT  8.680 4.000 10.600 4.240 ;
        RECT  10.360 4.000 10.600 4.530 ;
        RECT  12.900 4.230 14.140 4.470 ;
        RECT  10.360 4.290 13.140 4.530 ;
        RECT  14.070 2.140 14.670 2.540 ;
        RECT  14.070 1.610 14.310 3.510 ;
        RECT  11.140 1.610 11.540 2.010 ;
        RECT  11.300 1.610 11.540 4.050 ;
        RECT  11.140 3.250 11.540 4.050 ;
        RECT  14.750 3.590 15.150 3.990 ;
        RECT  12.400 3.750 15.150 3.990 ;
        RECT  14.910 1.610 15.150 3.990 ;
        RECT  11.140 3.810 12.700 4.050 ;
        RECT  16.120 1.860 17.110 2.100 ;
        RECT  16.870 2.360 17.500 2.600 ;
        RECT  16.870 1.860 17.110 3.530 ;
        RECT  16.050 3.290 17.110 3.530 ;
        RECT  5.390 1.130 18.500 1.370 ;
        RECT  18.220 1.130 18.500 3.510 ;
        RECT  11.960 1.130 12.200 3.570 ;
        RECT  5.390 1.130 5.630 3.650 ;
        RECT  5.170 3.250 5.630 3.650 ;
        RECT  17.480 1.720 17.980 2.120 ;
        RECT  17.350 3.290 17.980 3.530 ;
        RECT  17.740 1.720 17.980 4.060 ;
        RECT  17.740 3.820 18.760 4.060 ;
        RECT  19.660 1.450 20.060 1.850 ;
        RECT  19.720 1.450 19.960 3.510 ;
        RECT  19.600 3.110 20.020 3.510 ;
        RECT  18.880 3.110 19.280 3.510 ;
        RECT  19.000 1.450 19.240 3.990 ;
        RECT  21.590 2.580 21.830 3.990 ;
        RECT  19.000 3.750 21.830 3.990 ;
        RECT  20.200 2.100 22.630 2.340 ;
        RECT  21.080 2.100 21.320 3.510 ;
        RECT  22.390 1.640 22.630 3.720 ;
        RECT  15.390 3.840 15.790 4.370 ;
        RECT  23.870 3.910 25.440 4.150 ;
        RECT  18.930 4.230 24.110 4.470 ;
        RECT  15.390 4.130 17.460 4.370 ;
        RECT  23.870 1.640 24.110 4.470 ;
        RECT  17.220 4.300 19.100 4.540 ;
        RECT  25.200 3.910 25.440 4.620 ;
        RECT  23.130 1.160 24.590 1.400 ;
        RECT  24.350 1.160 24.590 1.940 ;
        RECT  24.350 1.700 26.200 1.940 ;
        RECT  25.960 1.840 26.540 2.090 ;
        RECT  23.130 1.160 23.370 3.720 ;
        RECT  25.880 1.220 27.020 1.460 ;
        RECT  26.780 1.220 27.020 2.570 ;
        RECT  26.780 2.170 27.270 2.570 ;
        RECT  26.050 2.330 27.270 2.570 ;
        RECT  24.870 3.270 26.290 3.510 ;
        RECT  26.050 2.330 26.290 3.670 ;
        RECT  25.890 3.270 26.290 3.670 ;
    END
END seprq1

MACRO sepfq4
    CLASS CORE ;
    FOREIGN sepfq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.515  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 2.220 8.900 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.340 1.800 5.780 2.040 ;
        RECT  4.540 1.460 4.980 2.040 ;
        RECT  4.340 1.800 4.580 2.510 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.882  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.300 2.460 ;
        RECT  2.530 2.020 3.300 2.420 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.886  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.490 1.350 21.370 1.750 ;
        RECT  20.970 1.020 21.370 1.750 ;
        RECT  20.670 2.020 21.220 2.460 ;
        RECT  19.030 3.060 21.070 3.460 ;
        RECT  20.670 1.350 21.070 3.460 ;
        RECT  20.330 3.060 20.730 3.900 ;
        RECT  19.490 1.020 19.890 1.750 ;
        RECT  19.030 3.060 19.430 3.960 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.533  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.290 2.260 0.690 2.660 ;
        RECT  0.120 2.020 0.500 2.460 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.370  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.270 2.020 7.780 2.460 ;
        RECT  7.270 2.020 7.670 2.970 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.380 2.090 13.940 2.480 ;
        RECT  13.500 2.020 13.940 2.480 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 21.840 5.600 ;
        RECT  20.930 4.220 21.330 5.600 ;
        RECT  19.590 4.260 19.990 5.600 ;
        RECT  18.510 2.900 18.750 5.600 ;
        RECT  16.560 4.620 16.960 5.600 ;
        RECT  13.680 4.340 14.080 5.600 ;
        RECT  12.490 4.210 12.730 5.600 ;
        RECT  8.870 4.480 9.270 5.600 ;
        RECT  6.430 4.170 6.830 5.600 ;
        RECT  2.860 3.960 3.260 5.600 ;
        RECT  0.750 3.560 1.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 21.840 0.740 ;
        RECT  20.230 0.000 20.630 1.110 ;
        RECT  18.750 0.000 19.150 1.170 ;
        RECT  17.460 0.000 17.860 1.050 ;
        RECT  13.550 0.000 13.790 1.200 ;
        RECT  9.520 0.000 9.920 0.890 ;
        RECT  7.040 0.000 7.280 1.200 ;
        RECT  3.030 0.000 3.270 1.200 ;
        RECT  0.150 0.000 0.550 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.170 1.780 ;
        RECT  0.930 2.330 1.510 2.570 ;
        RECT  0.930 1.540 1.170 3.320 ;
        RECT  0.230 3.080 1.170 3.320 ;
        RECT  0.230 3.080 0.470 4.620 ;
        RECT  1.530 1.430 2.040 1.830 ;
        RECT  1.800 2.170 2.250 2.570 ;
        RECT  1.800 1.430 2.040 3.280 ;
        RECT  1.490 3.040 2.040 3.280 ;
        RECT  2.210 0.980 2.770 1.220 ;
        RECT  2.530 0.980 2.770 1.680 ;
        RECT  2.530 1.440 3.780 1.680 ;
        RECT  6.140 1.840 6.380 2.530 ;
        RECT  4.990 2.290 6.380 2.530 ;
        RECT  3.540 1.440 3.780 3.450 ;
        RECT  4.990 2.290 5.230 3.450 ;
        RECT  2.280 3.210 5.230 3.450 ;
        RECT  2.280 3.210 2.520 3.700 ;
        RECT  2.200 3.460 2.440 4.360 ;
        RECT  8.690 1.740 9.380 1.980 ;
        RECT  9.140 2.600 9.950 2.840 ;
        RECT  9.140 1.740 9.380 3.500 ;
        RECT  8.300 3.260 9.380 3.500 ;
        RECT  10.090 1.780 11.020 2.020 ;
        RECT  10.090 1.700 10.490 2.100 ;
        RECT  10.190 1.700 10.430 3.370 ;
        RECT  9.620 3.130 10.430 3.370 ;
        RECT  7.600 0.980 8.560 1.220 ;
        RECT  5.050 0.980 6.800 1.220 ;
        RECT  10.160 0.980 11.500 1.220 ;
        RECT  8.160 1.140 10.400 1.380 ;
        RECT  6.560 0.980 6.800 1.680 ;
        RECT  7.600 0.980 7.840 1.680 ;
        RECT  6.560 1.440 7.840 1.680 ;
        RECT  11.260 0.980 11.500 2.500 ;
        RECT  10.670 2.260 11.500 2.500 ;
        RECT  6.790 1.440 7.030 3.450 ;
        RECT  5.470 3.210 7.920 3.450 ;
        RECT  7.680 3.210 7.920 3.760 ;
        RECT  5.470 3.210 5.710 3.940 ;
        RECT  4.530 3.690 5.710 3.940 ;
        RECT  10.670 2.260 10.910 4.140 ;
        RECT  10.140 3.900 10.910 4.140 ;
        RECT  12.230 1.460 12.820 1.700 ;
        RECT  12.230 1.460 12.470 3.460 ;
        RECT  11.810 3.220 12.470 3.460 ;
        RECT  11.740 0.980 13.310 1.220 ;
        RECT  13.070 0.980 13.310 1.780 ;
        RECT  13.070 1.540 14.480 1.780 ;
        RECT  14.240 1.540 14.480 2.480 ;
        RECT  11.740 0.980 11.980 2.980 ;
        RECT  11.150 2.740 11.980 2.980 ;
        RECT  11.150 2.740 11.390 3.510 ;
        RECT  14.670 0.990 15.070 1.390 ;
        RECT  12.710 2.010 12.950 3.040 ;
        RECT  14.720 0.990 14.960 3.040 ;
        RECT  12.710 2.800 14.960 3.040 ;
        RECT  13.190 3.860 14.560 4.100 ;
        RECT  14.320 4.050 17.440 4.290 ;
        RECT  13.190 3.860 13.430 4.580 ;
        RECT  12.970 4.180 13.430 4.580 ;
        RECT  17.200 4.050 17.440 4.620 ;
        RECT  16.180 1.460 16.740 1.700 ;
        RECT  16.500 2.800 17.560 3.040 ;
        RECT  12.710 3.380 14.960 3.620 ;
        RECT  16.500 1.460 16.740 3.650 ;
        RECT  14.720 3.410 16.740 3.650 ;
        RECT  5.950 3.690 7.320 3.930 ;
        RECT  12.710 3.380 12.950 3.940 ;
        RECT  11.930 3.700 12.950 3.940 ;
        RECT  7.080 3.690 7.320 4.240 ;
        RECT  7.080 4.000 9.750 4.240 ;
        RECT  9.510 4.000 9.750 4.620 ;
        RECT  5.950 3.690 6.190 4.500 ;
        RECT  4.900 4.260 6.190 4.500 ;
        RECT  11.930 3.700 12.170 4.620 ;
        RECT  9.510 4.380 12.170 4.620 ;
        RECT  15.490 0.980 17.220 1.220 ;
        RECT  15.490 0.980 15.730 1.860 ;
        RECT  15.200 1.620 15.730 1.860 ;
        RECT  16.980 0.980 17.220 2.180 ;
        RECT  16.980 1.940 18.300 2.180 ;
        RECT  15.200 1.620 15.440 3.140 ;
        RECT  17.990 1.410 19.100 1.650 ;
        RECT  18.860 2.010 20.430 2.410 ;
        RECT  18.860 1.410 19.100 2.660 ;
        RECT  18.030 2.420 19.100 2.660 ;
        RECT  18.030 2.420 18.270 4.620 ;
        RECT  17.690 4.380 18.270 4.620 ;
    END
END sepfq4

MACRO sepfq2
    CLASS CORE ;
    FOREIGN sepfq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.515  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 2.220 8.900 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.340 1.800 5.780 2.040 ;
        RECT  4.540 1.460 4.980 2.040 ;
        RECT  4.340 1.800 4.580 2.510 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.882  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.300 2.460 ;
        RECT  2.530 2.020 3.300 2.420 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.040 2.690 20.040 3.020 ;
        RECT  19.660 1.380 20.040 3.020 ;
        RECT  19.250 1.380 20.040 1.780 ;
        RECT  19.040 2.690 19.440 4.330 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.533  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.290 2.260 0.690 2.660 ;
        RECT  0.120 2.020 0.500 2.460 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.370  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.270 2.020 7.780 2.460 ;
        RECT  7.270 2.020 7.670 2.970 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.380 2.080 13.940 2.480 ;
        RECT  13.500 2.020 13.940 2.480 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.160 5.600 ;
        RECT  19.690 3.260 19.930 5.600 ;
        RECT  18.480 4.620 18.880 5.600 ;
        RECT  16.520 4.620 16.920 5.600 ;
        RECT  13.680 4.340 14.080 5.600 ;
        RECT  12.490 4.210 12.730 5.600 ;
        RECT  8.870 4.480 9.270 5.600 ;
        RECT  6.510 4.170 6.750 5.600 ;
        RECT  2.860 3.960 3.260 5.600 ;
        RECT  0.750 3.580 1.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.160 0.740 ;
        RECT  18.680 0.000 19.080 0.990 ;
        RECT  13.550 0.000 13.790 1.300 ;
        RECT  9.520 0.000 9.920 0.890 ;
        RECT  7.040 0.000 7.280 1.200 ;
        RECT  3.030 0.000 3.270 1.200 ;
        RECT  0.150 0.000 0.550 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.170 1.780 ;
        RECT  0.930 2.250 1.510 2.650 ;
        RECT  0.930 1.540 1.170 3.340 ;
        RECT  0.230 3.100 1.170 3.340 ;
        RECT  0.230 3.100 0.470 4.620 ;
        RECT  1.530 1.430 2.040 1.830 ;
        RECT  1.800 2.170 2.250 2.570 ;
        RECT  1.800 1.430 2.040 3.280 ;
        RECT  1.490 3.040 2.040 3.280 ;
        RECT  2.210 0.980 2.770 1.220 ;
        RECT  2.530 0.980 2.770 1.680 ;
        RECT  2.530 1.440 3.780 1.680 ;
        RECT  6.140 1.840 6.380 2.530 ;
        RECT  5.010 2.290 6.380 2.530 ;
        RECT  3.540 1.440 3.780 3.450 ;
        RECT  5.010 2.290 5.250 3.450 ;
        RECT  2.280 3.210 5.250 3.450 ;
        RECT  2.280 3.210 2.520 3.700 ;
        RECT  2.200 3.460 2.440 4.360 ;
        RECT  8.690 1.740 9.380 1.980 ;
        RECT  9.140 2.600 9.950 2.840 ;
        RECT  9.140 1.740 9.380 3.500 ;
        RECT  8.300 3.260 9.380 3.500 ;
        RECT  10.090 1.780 11.020 2.020 ;
        RECT  10.090 1.700 10.490 2.100 ;
        RECT  10.190 1.700 10.430 3.370 ;
        RECT  9.620 3.130 10.430 3.370 ;
        RECT  5.050 0.980 6.800 1.220 ;
        RECT  7.600 0.980 8.560 1.220 ;
        RECT  10.160 0.980 11.500 1.220 ;
        RECT  6.560 0.980 6.800 1.680 ;
        RECT  8.160 1.220 10.400 1.460 ;
        RECT  7.600 0.980 7.840 1.680 ;
        RECT  6.560 1.440 7.840 1.680 ;
        RECT  11.260 0.980 11.500 2.500 ;
        RECT  10.670 2.260 11.500 2.500 ;
        RECT  6.790 1.440 7.030 3.450 ;
        RECT  5.490 3.210 7.920 3.450 ;
        RECT  7.680 3.210 7.920 3.760 ;
        RECT  5.490 3.210 5.730 3.940 ;
        RECT  4.530 3.700 5.730 3.940 ;
        RECT  10.670 2.260 10.910 4.140 ;
        RECT  10.140 3.900 10.910 4.140 ;
        RECT  12.230 1.460 12.820 1.700 ;
        RECT  12.230 1.460 12.470 3.460 ;
        RECT  11.810 3.220 12.470 3.460 ;
        RECT  11.740 0.980 13.310 1.220 ;
        RECT  13.070 0.980 13.310 1.780 ;
        RECT  13.070 1.540 14.480 1.780 ;
        RECT  14.240 1.540 14.480 2.480 ;
        RECT  11.740 0.980 11.980 2.980 ;
        RECT  11.150 2.740 11.980 2.980 ;
        RECT  11.150 2.740 11.390 3.510 ;
        RECT  14.670 0.980 15.070 1.380 ;
        RECT  12.710 2.010 12.950 3.040 ;
        RECT  14.720 0.980 14.960 3.040 ;
        RECT  12.710 2.800 14.960 3.040 ;
        RECT  13.190 3.860 14.560 4.100 ;
        RECT  14.320 4.050 17.400 4.290 ;
        RECT  13.190 3.860 13.430 4.580 ;
        RECT  12.970 4.180 13.430 4.580 ;
        RECT  17.160 4.050 17.400 4.620 ;
        RECT  16.180 1.460 16.740 1.700 ;
        RECT  16.500 2.800 17.560 3.040 ;
        RECT  12.710 3.380 14.960 3.620 ;
        RECT  16.500 1.460 16.740 3.650 ;
        RECT  14.720 3.410 16.740 3.650 ;
        RECT  5.970 3.690 7.320 3.930 ;
        RECT  12.710 3.380 12.950 3.940 ;
        RECT  11.930 3.700 12.950 3.940 ;
        RECT  7.080 3.690 7.320 4.240 ;
        RECT  7.080 4.000 9.750 4.240 ;
        RECT  9.510 4.000 9.750 4.620 ;
        RECT  5.970 3.690 6.210 4.500 ;
        RECT  4.900 4.260 6.210 4.500 ;
        RECT  11.930 3.700 12.170 4.620 ;
        RECT  9.510 4.380 12.170 4.620 ;
        RECT  15.490 0.980 17.220 1.220 ;
        RECT  15.490 0.980 15.730 1.860 ;
        RECT  15.200 1.620 15.730 1.860 ;
        RECT  16.980 0.980 17.220 2.250 ;
        RECT  16.980 2.010 18.250 2.250 ;
        RECT  15.200 1.620 15.440 3.140 ;
        RECT  17.910 1.480 18.730 1.720 ;
        RECT  18.490 2.050 19.270 2.450 ;
        RECT  18.490 1.480 18.730 2.730 ;
        RECT  18.000 2.490 18.730 2.730 ;
        RECT  18.000 2.490 18.240 4.620 ;
        RECT  17.690 4.380 18.240 4.620 ;
    END
END sepfq2

MACRO sepfq1
    CLASS CORE ;
    FOREIGN sepfq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.515  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.820 2.200 9.220 2.600 ;
        RECT  8.460 2.580 9.060 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.490 1.600 5.890 2.000 ;
        RECT  4.370 2.250 5.810 2.490 ;
        RECT  5.570 1.600 5.810 2.490 ;
        RECT  4.370 2.170 4.980 2.490 ;
        RECT  4.540 2.020 4.980 2.490 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.898  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.600 2.020 3.300 2.460 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.069  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  20.780 2.020 21.160 2.460 ;
        RECT  20.790 1.620 21.030 3.470 ;
        RECT  20.740 1.060 20.980 1.860 ;
        RECT  20.780 1.620 21.030 2.460 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.529  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.290 2.260 0.690 2.820 ;
        RECT  0.120 2.580 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.370  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.580 7.710 2.840 ;
        RECT  7.310 2.440 7.710 2.840 ;
        RECT  6.780 2.580 7.220 3.020 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.860 2.020 14.500 2.500 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 21.280 5.600 ;
        RECT  19.980 3.970 20.380 5.600 ;
        RECT  18.020 4.550 18.420 5.600 ;
        RECT  15.710 4.380 15.950 5.600 ;
        RECT  15.400 4.380 15.950 4.620 ;
        RECT  13.330 4.300 13.570 5.600 ;
        RECT  9.280 4.480 9.680 5.600 ;
        RECT  6.770 4.340 7.180 5.600 ;
        RECT  2.850 3.690 3.250 5.600 ;
        RECT  0.750 4.030 1.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 21.280 0.740 ;
        RECT  19.890 0.000 20.290 0.980 ;
        RECT  18.470 0.000 18.710 1.380 ;
        RECT  13.620 0.000 14.020 1.290 ;
        RECT  9.560 0.000 9.960 0.900 ;
        RECT  6.880 0.000 7.280 1.250 ;
        RECT  2.980 0.000 3.380 0.970 ;
        RECT  0.740 0.000 1.140 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.770 1.170 2.010 ;
        RECT  0.930 2.330 1.490 2.570 ;
        RECT  0.930 1.770 1.170 3.670 ;
        RECT  0.150 3.430 1.170 3.670 ;
        RECT  1.590 1.310 1.830 2.060 ;
        RECT  1.590 1.820 2.090 2.060 ;
        RECT  1.850 1.820 2.090 3.430 ;
        RECT  1.470 3.190 2.090 3.430 ;
        RECT  2.210 1.180 2.760 1.420 ;
        RECT  2.520 1.210 4.090 1.450 ;
        RECT  3.850 1.210 4.090 2.970 ;
        RECT  3.050 2.730 6.490 2.970 ;
        RECT  6.250 2.040 6.490 2.970 ;
        RECT  2.360 2.800 3.290 3.040 ;
        RECT  2.360 2.800 2.600 3.350 ;
        RECT  8.790 1.710 9.770 1.950 ;
        RECT  9.530 2.520 10.090 2.920 ;
        RECT  9.530 1.710 9.770 3.500 ;
        RECT  8.710 3.260 9.770 3.500 ;
        RECT  10.330 1.630 10.730 2.120 ;
        RECT  10.330 1.880 11.170 2.120 ;
        RECT  10.930 1.880 11.170 2.470 ;
        RECT  10.330 1.630 10.570 3.430 ;
        RECT  10.010 3.190 10.570 3.430 ;
        RECT  4.970 0.980 6.480 1.220 ;
        RECT  8.080 1.150 11.650 1.390 ;
        RECT  6.240 0.980 6.480 1.730 ;
        RECT  8.080 1.140 8.480 1.540 ;
        RECT  11.030 1.150 11.650 1.550 ;
        RECT  6.240 1.490 8.400 1.730 ;
        RECT  11.410 1.150 11.650 2.950 ;
        RECT  11.030 2.710 11.650 2.950 ;
        RECT  4.590 3.250 6.360 3.490 ;
        RECT  7.450 3.250 8.300 3.490 ;
        RECT  7.950 1.490 8.190 3.490 ;
        RECT  6.120 3.310 7.690 3.550 ;
        RECT  8.060 3.250 8.300 3.910 ;
        RECT  11.030 2.710 11.270 4.140 ;
        RECT  10.720 3.900 11.270 4.140 ;
        RECT  12.370 3.190 13.090 3.430 ;
        RECT  12.630 1.660 12.870 3.430 ;
        RECT  12.850 3.220 14.120 3.460 ;
        RECT  12.370 3.190 12.610 3.740 ;
        RECT  11.890 0.980 13.350 1.220 ;
        RECT  14.260 0.980 15.780 1.220 ;
        RECT  13.110 0.980 13.350 1.780 ;
        RECT  14.260 0.980 14.500 1.780 ;
        RECT  13.110 1.540 14.500 1.780 ;
        RECT  15.540 0.980 15.780 2.700 ;
        RECT  15.350 2.300 15.780 2.700 ;
        RECT  11.890 0.980 12.130 3.430 ;
        RECT  11.540 3.190 12.130 3.430 ;
        RECT  11.540 3.190 11.780 3.740 ;
        RECT  14.740 1.640 15.300 1.880 ;
        RECT  14.740 1.640 14.980 3.180 ;
        RECT  13.110 2.470 13.510 2.870 ;
        RECT  13.270 2.740 14.980 2.980 ;
        RECT  14.420 2.940 16.120 3.180 ;
        RECT  17.190 1.460 17.740 1.700 ;
        RECT  17.500 1.460 17.740 2.950 ;
        RECT  17.340 2.710 17.580 3.710 ;
        RECT  14.440 3.420 17.070 3.660 ;
        RECT  18.790 3.140 19.040 3.710 ;
        RECT  16.830 3.470 19.040 3.710 ;
        RECT  14.440 3.420 14.680 3.940 ;
        RECT  12.850 3.700 14.680 3.940 ;
        RECT  6.050 3.860 7.710 4.100 ;
        RECT  8.790 3.980 10.160 4.220 ;
        RECT  5.130 4.020 6.290 4.260 ;
        RECT  7.470 3.860 7.710 4.620 ;
        RECT  9.920 3.980 10.160 4.620 ;
        RECT  5.130 4.020 5.370 4.580 ;
        RECT  8.790 3.980 9.030 4.620 ;
        RECT  7.470 4.380 9.030 4.620 ;
        RECT  12.850 3.700 13.090 4.620 ;
        RECT  9.920 4.380 13.090 4.620 ;
        RECT  14.920 3.900 16.560 4.140 ;
        RECT  16.300 3.950 18.900 4.190 ;
        RECT  18.660 3.950 18.900 4.620 ;
        RECT  14.920 3.900 15.160 4.500 ;
        RECT  13.870 4.260 15.160 4.500 ;
        RECT  18.660 4.380 19.210 4.620 ;
        RECT  16.670 0.980 18.220 1.220 ;
        RECT  16.250 1.250 16.910 1.490 ;
        RECT  17.980 0.980 18.220 1.950 ;
        RECT  17.980 1.710 19.150 1.950 ;
        RECT  18.910 1.710 19.150 2.420 ;
        RECT  16.670 0.980 16.910 2.310 ;
        RECT  18.910 2.020 19.320 2.420 ;
        RECT  16.770 2.070 17.010 3.180 ;
        RECT  16.460 2.940 17.010 3.180 ;
        RECT  19.120 1.110 19.680 1.350 ;
        RECT  19.440 1.220 20.040 1.460 ;
        RECT  19.800 2.040 20.200 2.440 ;
        RECT  19.800 1.220 20.040 3.160 ;
        RECT  19.490 2.920 20.040 3.160 ;
        RECT  19.490 2.920 19.730 3.470 ;
    END
END sepfq1

MACRO senrq4
    CLASS CORE ;
    FOREIGN senrq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 2.020 8.900 2.460 ;
        RECT  8.350 2.200 8.750 2.600 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 4.980 2.460 ;
        RECT  4.140 2.040 4.980 2.440 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.880 2.510 6.320 2.910 ;
        RECT  5.880 1.970 6.120 2.910 ;
        RECT  5.220 1.970 6.120 2.210 ;
        RECT  5.220 1.540 5.460 2.210 ;
        RECT  4.020 1.540 5.460 1.780 ;
        RECT  3.060 1.460 4.260 1.700 ;
        RECT  3.060 1.460 3.300 2.460 ;
        RECT  2.760 2.220 3.160 2.810 ;
        RECT  2.860 2.020 3.300 2.460 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.074  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.100 3.100 19.480 3.610 ;
        RECT  19.050 1.260 19.450 1.660 ;
        RECT  16.810 3.930 19.340 4.170 ;
        RECT  19.100 1.260 19.340 4.170 ;
        RECT  17.680 1.340 19.450 1.580 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.449  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.710 0.540 3.110 ;
        RECT  0.120 2.020 0.500 2.880 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.387  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.020 7.780 2.460 ;
        RECT  7.170 2.030 7.780 2.430 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.600 5.600 ;
        RECT  19.050 4.620 19.450 5.600 ;
        RECT  17.750 4.620 18.150 5.600 ;
        RECT  16.440 4.620 16.840 5.600 ;
        RECT  15.170 4.620 15.570 5.600 ;
        RECT  12.290 4.710 12.690 5.600 ;
        RECT  8.920 4.710 9.320 5.600 ;
        RECT  6.180 4.620 6.580 5.600 ;
        RECT  2.950 4.370 3.190 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.600 0.740 ;
        RECT  18.240 0.000 18.640 0.980 ;
        RECT  16.910 0.000 17.310 0.890 ;
        RECT  15.640 0.000 16.040 0.980 ;
        RECT  12.590 0.000 12.990 0.890 ;
        RECT  9.050 0.000 9.450 0.890 ;
        RECT  6.280 0.000 6.680 1.200 ;
        RECT  2.410 0.000 2.830 0.930 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.420 0.980 1.660 ;
        RECT  0.740 1.420 0.980 2.240 ;
        RECT  0.740 2.000 1.260 2.240 ;
        RECT  1.020 2.000 1.260 3.690 ;
        RECT  0.150 3.450 1.260 3.690 ;
        RECT  1.220 0.980 1.940 1.220 ;
        RECT  1.220 0.980 1.460 1.710 ;
        RECT  1.220 1.470 1.740 1.710 ;
        RECT  1.500 1.470 1.740 2.490 ;
        RECT  1.500 2.250 2.030 2.490 ;
        RECT  1.790 2.250 2.030 2.980 ;
        RECT  1.570 2.740 1.810 3.680 ;
        RECT  2.060 1.590 2.520 1.990 ;
        RECT  3.540 2.180 3.780 3.360 ;
        RECT  2.280 3.120 3.780 3.360 ;
        RECT  2.280 1.590 2.520 3.620 ;
        RECT  2.200 3.380 2.440 4.480 ;
        RECT  8.280 1.540 9.380 1.780 ;
        RECT  9.140 1.540 9.380 2.670 ;
        RECT  9.140 2.180 9.620 2.600 ;
        RECT  9.120 2.560 9.440 2.670 ;
        RECT  9.120 2.560 9.360 3.210 ;
        RECT  8.230 2.970 9.360 3.210 ;
        RECT  9.720 1.300 9.960 1.940 ;
        RECT  9.720 1.700 10.220 1.940 ;
        RECT  9.980 1.700 10.220 3.180 ;
        RECT  9.610 2.940 10.220 3.180 ;
        RECT  9.610 2.940 9.850 3.510 ;
        RECT  4.330 0.980 5.390 1.220 ;
        RECT  5.170 1.060 5.940 1.300 ;
        RECT  10.340 0.980 10.740 1.380 ;
        RECT  6.920 1.170 7.880 1.410 ;
        RECT  5.700 1.060 5.940 1.730 ;
        RECT  6.920 1.170 7.160 1.730 ;
        RECT  5.700 1.490 7.160 1.730 ;
        RECT  6.560 1.490 6.800 3.700 ;
        RECT  5.020 3.460 7.990 3.700 ;
        RECT  4.540 3.560 5.260 3.800 ;
        RECT  7.750 3.560 8.920 3.800 ;
        RECT  8.680 3.750 10.740 3.990 ;
        RECT  10.500 0.980 10.740 4.070 ;
        RECT  10.230 3.670 10.740 4.070 ;
        RECT  11.670 1.650 12.220 1.890 ;
        RECT  11.670 1.650 11.910 2.150 ;
        RECT  11.540 1.910 11.780 3.570 ;
        RECT  11.670 3.330 11.910 3.970 ;
        RECT  10.980 1.130 12.830 1.410 ;
        RECT  10.980 1.130 11.480 1.500 ;
        RECT  10.980 1.130 11.400 1.600 ;
        RECT  12.590 1.130 12.830 2.150 ;
        RECT  12.830 1.900 13.070 2.500 ;
        RECT  10.980 1.130 11.220 3.400 ;
        RECT  13.310 1.070 13.760 1.470 ;
        RECT  13.310 1.070 13.550 3.080 ;
        RECT  12.020 2.470 12.260 3.090 ;
        RECT  13.260 2.820 13.500 3.360 ;
        RECT  12.730 3.120 13.500 3.360 ;
        RECT  12.150 2.850 12.390 3.640 ;
        RECT  12.150 3.400 12.970 3.640 ;
        RECT  12.730 3.120 12.970 3.980 ;
        RECT  12.730 3.740 13.290 3.980 ;
        RECT  13.830 1.840 14.070 2.770 ;
        RECT  13.900 2.510 14.140 3.360 ;
        RECT  5.240 2.460 5.640 2.860 ;
        RECT  4.030 2.720 5.450 2.960 ;
        RECT  4.030 2.720 4.520 3.120 ;
        RECT  4.030 2.720 4.270 4.280 ;
        RECT  4.030 4.040 8.440 4.280 ;
        RECT  14.950 1.620 15.190 4.320 ;
        RECT  14.370 4.080 15.190 4.320 ;
        RECT  8.200 4.230 9.980 4.470 ;
        RECT  10.980 4.230 13.200 4.470 ;
        RECT  9.740 4.320 11.220 4.560 ;
        RECT  14.370 4.080 14.770 4.620 ;
        RECT  12.960 4.380 14.770 4.620 ;
        RECT  14.100 1.170 15.410 1.380 ;
        RECT  14.100 1.180 15.430 1.380 ;
        RECT  14.100 1.190 15.470 1.380 ;
        RECT  14.100 1.210 15.500 1.380 ;
        RECT  14.100 1.140 15.330 1.380 ;
        RECT  15.260 1.220 16.250 1.390 ;
        RECT  15.290 1.220 16.250 1.400 ;
        RECT  15.310 1.220 16.250 1.410 ;
        RECT  15.330 1.150 15.360 1.420 ;
        RECT  15.340 1.220 16.250 1.430 ;
        RECT  15.350 1.220 16.250 1.440 ;
        RECT  15.360 1.160 15.390 1.450 ;
        RECT  15.370 1.220 16.250 1.460 ;
        RECT  14.100 1.070 14.670 1.470 ;
        RECT  16.010 1.220 16.250 2.770 ;
        RECT  13.820 3.600 14.670 3.840 ;
        RECT  14.430 1.070 14.670 3.840 ;
        RECT  13.630 3.660 14.060 4.060 ;
        RECT  16.490 2.260 18.860 2.660 ;
        RECT  15.490 1.700 15.730 3.360 ;
        RECT  16.490 1.300 16.730 3.360 ;
        RECT  15.490 3.120 16.730 3.360 ;
    END
END senrq4

MACRO senrq2
    CLASS CORE ;
    FOREIGN senrq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.320 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.580 16.360 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.940 2.250 13.380 3.020 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.397  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.700 2.580 7.310 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  25.130 3.150 25.630 4.140 ;
        RECT  25.390 1.460 25.630 4.140 ;
        RECT  25.170 1.460 25.630 1.880 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.020 0.980 2.900 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.280 1.640 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 26.320 5.600 ;
        RECT  25.700 4.450 26.100 5.600 ;
        RECT  24.390 4.450 24.790 5.600 ;
        RECT  23.200 3.120 23.440 5.600 ;
        RECT  20.230 4.670 20.630 5.600 ;
        RECT  16.310 4.640 16.710 5.600 ;
        RECT  14.640 4.710 15.040 5.600 ;
        RECT  13.390 4.710 13.790 5.600 ;
        RECT  9.670 4.480 10.070 5.600 ;
        RECT  8.200 3.770 8.440 5.600 ;
        RECT  6.900 3.770 7.140 5.600 ;
        RECT  6.000 3.850 6.240 5.600 ;
        RECT  3.930 4.090 4.170 5.600 ;
        RECT  1.660 4.460 2.060 5.600 ;
        RECT  0.970 3.290 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 26.320 0.740 ;
        RECT  25.740 0.000 26.140 1.140 ;
        RECT  24.430 0.000 24.830 1.140 ;
        RECT  23.240 0.000 23.480 1.850 ;
        RECT  20.040 0.000 20.280 1.800 ;
        RECT  16.460 0.000 16.860 0.890 ;
        RECT  15.050 0.000 15.450 0.890 ;
        RECT  13.070 0.000 13.470 0.890 ;
        RECT  10.170 0.000 10.570 0.890 ;
        RECT  8.130 0.000 8.530 0.890 ;
        RECT  6.180 0.000 6.600 0.890 ;
        RECT  4.190 0.000 4.430 1.470 ;
        RECT  1.660 0.000 2.060 1.140 ;
        RECT  0.760 0.000 1.180 1.180 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 1.520 0.470 1.920 ;
        RECT  0.220 1.520 0.460 4.620 ;
        RECT  0.220 3.290 0.470 4.620 ;
        RECT  1.570 1.530 2.120 1.930 ;
        RECT  1.880 2.270 2.990 2.510 ;
        RECT  1.880 1.530 2.120 3.650 ;
        RECT  1.630 3.260 2.120 3.650 ;
        RECT  2.430 0.980 2.990 1.380 ;
        RECT  2.670 0.980 2.990 1.910 ;
        RECT  2.670 1.630 3.470 1.910 ;
        RECT  3.230 1.630 3.470 2.990 ;
        RECT  2.480 2.750 3.470 2.990 ;
        RECT  2.480 2.750 2.720 4.620 ;
        RECT  2.430 4.220 2.830 4.620 ;
        RECT  3.230 1.150 3.950 1.390 ;
        RECT  3.710 2.800 4.450 3.040 ;
        RECT  3.710 1.150 3.950 3.610 ;
        RECT  2.960 3.370 3.950 3.610 ;
        RECT  2.960 3.370 3.360 3.770 ;
        RECT  4.570 1.830 4.930 2.230 ;
        RECT  4.690 1.830 4.930 3.750 ;
        RECT  4.430 3.350 4.930 3.750 ;
        RECT  6.000 1.610 6.580 1.850 ;
        RECT  6.000 1.610 6.240 3.510 ;
        RECT  9.440 1.610 9.680 2.500 ;
        RECT  9.160 2.260 10.280 2.500 ;
        RECT  9.160 2.260 9.400 3.740 ;
        RECT  10.170 1.690 10.760 1.930 ;
        RECT  10.520 1.690 10.760 3.740 ;
        RECT  10.520 2.510 11.050 2.910 ;
        RECT  10.520 2.510 10.840 3.740 ;
        RECT  10.440 3.340 10.840 3.740 ;
        RECT  12.460 1.610 12.880 2.010 ;
        RECT  12.460 1.610 12.700 3.510 ;
        RECT  12.460 3.270 13.020 3.510 ;
        RECT  6.900 1.620 7.860 1.860 ;
        RECT  7.620 1.620 7.860 3.510 ;
        RECT  7.540 3.110 7.940 3.510 ;
        RECT  7.540 3.270 8.920 3.510 ;
        RECT  8.680 3.270 8.920 4.240 ;
        RECT  8.680 4.000 10.600 4.240 ;
        RECT  10.360 4.000 10.600 4.530 ;
        RECT  12.900 4.230 14.140 4.470 ;
        RECT  10.360 4.290 13.140 4.530 ;
        RECT  13.930 1.610 14.170 2.540 ;
        RECT  13.930 2.140 14.530 2.540 ;
        RECT  14.070 2.140 14.310 3.510 ;
        RECT  11.000 1.610 11.540 2.010 ;
        RECT  14.790 1.630 15.450 2.030 ;
        RECT  11.300 1.610 11.540 4.050 ;
        RECT  11.140 3.250 11.540 4.050 ;
        RECT  12.400 3.750 15.030 3.990 ;
        RECT  11.140 3.810 12.700 4.050 ;
        RECT  14.790 1.630 15.030 4.350 ;
        RECT  15.850 1.860 16.840 2.100 ;
        RECT  16.600 2.440 17.230 2.680 ;
        RECT  16.600 1.860 16.840 3.530 ;
        RECT  15.780 3.290 16.840 3.530 ;
        RECT  5.390 1.130 18.230 1.370 ;
        RECT  17.710 0.980 18.230 1.400 ;
        RECT  11.820 1.130 12.060 2.900 ;
        RECT  17.990 0.980 18.230 3.470 ;
        RECT  11.960 2.600 12.200 3.570 ;
        RECT  5.390 1.130 5.630 3.650 ;
        RECT  5.170 3.250 5.630 3.650 ;
        RECT  17.180 1.780 17.710 2.180 ;
        RECT  17.080 3.290 17.710 3.530 ;
        RECT  17.470 1.780 17.710 4.020 ;
        RECT  17.470 3.780 18.490 4.020 ;
        RECT  19.230 1.450 19.540 3.470 ;
        RECT  19.230 3.070 19.790 3.470 ;
        RECT  18.560 1.450 18.800 2.700 ;
        RECT  20.030 2.620 20.860 2.860 ;
        RECT  18.730 2.400 18.970 3.950 ;
        RECT  20.030 2.620 20.270 3.950 ;
        RECT  18.730 3.710 20.270 3.950 ;
        RECT  20.790 1.450 21.030 2.300 ;
        RECT  19.780 2.060 21.390 2.300 ;
        RECT  21.150 2.060 21.390 3.390 ;
        RECT  20.820 3.150 21.390 3.390 ;
        RECT  22.280 1.480 22.520 3.950 ;
        RECT  22.280 3.160 22.760 3.950 ;
        RECT  20.510 3.710 22.760 3.950 ;
        RECT  15.270 3.420 15.510 4.370 ;
        RECT  18.660 4.190 20.750 4.430 ;
        RECT  15.270 4.130 17.250 4.370 ;
        RECT  20.510 3.710 20.750 4.430 ;
        RECT  17.010 4.300 18.900 4.540 ;
        RECT  21.520 1.000 23.000 1.240 ;
        RECT  21.520 1.000 21.930 1.850 ;
        RECT  22.760 1.000 23.000 2.380 ;
        RECT  22.760 2.140 23.970 2.380 ;
        RECT  21.690 1.000 21.930 3.470 ;
        RECT  23.860 1.610 24.450 1.850 ;
        RECT  24.210 1.610 24.450 2.860 ;
        RECT  24.210 2.610 25.150 2.860 ;
        RECT  22.760 2.620 25.150 2.860 ;
        RECT  23.900 2.620 24.140 3.470 ;
    END
END senrq2

MACRO senrq1
    CLASS CORE ;
    FOREIGN senrq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.760 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.580 16.360 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.940 2.250 13.380 3.020 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.397  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.700 2.580 7.310 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  25.160 3.150 25.630 4.140 ;
        RECT  25.390 1.460 25.630 4.140 ;
        RECT  25.210 1.460 25.630 1.880 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.020 0.980 2.900 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.280 1.640 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 25.760 5.600 ;
        RECT  24.390 4.450 24.790 5.600 ;
        RECT  23.200 3.120 23.440 5.600 ;
        RECT  20.230 4.670 20.630 5.600 ;
        RECT  16.310 4.640 16.710 5.600 ;
        RECT  14.640 4.710 15.040 5.600 ;
        RECT  13.390 4.710 13.790 5.600 ;
        RECT  9.670 4.480 10.070 5.600 ;
        RECT  8.200 3.770 8.440 5.600 ;
        RECT  6.900 3.770 7.140 5.600 ;
        RECT  6.000 3.850 6.240 5.600 ;
        RECT  3.930 4.090 4.170 5.600 ;
        RECT  1.660 4.460 2.060 5.600 ;
        RECT  0.970 3.290 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 25.760 0.740 ;
        RECT  24.470 0.000 24.870 1.140 ;
        RECT  23.240 0.000 23.480 1.850 ;
        RECT  20.040 0.000 20.280 1.800 ;
        RECT  16.460 0.000 16.860 0.890 ;
        RECT  15.050 0.000 15.450 0.890 ;
        RECT  13.070 0.000 13.470 0.890 ;
        RECT  10.170 0.000 10.570 0.890 ;
        RECT  8.130 0.000 8.530 0.890 ;
        RECT  6.180 0.000 6.600 0.890 ;
        RECT  4.190 0.000 4.430 1.470 ;
        RECT  1.660 0.000 2.060 1.140 ;
        RECT  0.760 0.000 1.180 1.180 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 1.520 0.470 1.920 ;
        RECT  0.220 1.520 0.460 4.620 ;
        RECT  0.220 3.290 0.470 4.620 ;
        RECT  1.570 1.530 2.120 1.930 ;
        RECT  1.880 2.270 2.990 2.510 ;
        RECT  1.880 1.530 2.120 3.650 ;
        RECT  1.630 3.260 2.120 3.650 ;
        RECT  2.430 0.980 2.990 1.380 ;
        RECT  2.670 0.980 2.990 1.910 ;
        RECT  2.670 1.630 3.470 1.910 ;
        RECT  3.230 1.630 3.470 2.990 ;
        RECT  2.480 2.750 3.470 2.990 ;
        RECT  2.480 2.750 2.720 4.620 ;
        RECT  2.430 4.220 2.830 4.620 ;
        RECT  3.230 1.150 3.950 1.390 ;
        RECT  3.710 2.800 4.450 3.040 ;
        RECT  3.710 1.150 3.950 3.610 ;
        RECT  2.960 3.370 3.950 3.610 ;
        RECT  2.960 3.370 3.360 3.770 ;
        RECT  4.570 1.830 4.930 2.230 ;
        RECT  4.690 1.830 4.930 3.750 ;
        RECT  4.430 3.350 4.930 3.750 ;
        RECT  6.000 1.610 6.580 1.850 ;
        RECT  6.000 1.610 6.240 3.510 ;
        RECT  9.440 1.610 9.680 2.500 ;
        RECT  9.160 2.260 10.280 2.500 ;
        RECT  9.160 2.260 9.400 3.740 ;
        RECT  10.170 1.690 10.760 1.930 ;
        RECT  10.520 1.690 10.760 3.740 ;
        RECT  10.520 2.510 11.050 2.910 ;
        RECT  10.520 2.510 10.840 3.740 ;
        RECT  10.440 3.340 10.840 3.740 ;
        RECT  12.460 1.610 12.880 2.010 ;
        RECT  12.460 1.610 12.700 3.510 ;
        RECT  12.460 3.270 13.020 3.510 ;
        RECT  6.900 1.620 7.860 1.860 ;
        RECT  7.620 1.620 7.860 3.510 ;
        RECT  7.540 3.110 7.940 3.510 ;
        RECT  7.540 3.270 8.920 3.510 ;
        RECT  8.680 3.270 8.920 4.240 ;
        RECT  8.680 4.000 10.600 4.240 ;
        RECT  10.360 4.000 10.600 4.530 ;
        RECT  12.900 4.230 14.140 4.470 ;
        RECT  10.360 4.290 13.140 4.530 ;
        RECT  13.930 1.610 14.170 2.540 ;
        RECT  13.930 2.140 14.530 2.540 ;
        RECT  14.070 2.140 14.310 3.510 ;
        RECT  11.000 1.610 11.540 2.010 ;
        RECT  14.790 1.630 15.450 2.030 ;
        RECT  11.300 1.610 11.540 4.050 ;
        RECT  11.140 3.250 11.540 4.050 ;
        RECT  12.400 3.750 15.030 3.990 ;
        RECT  11.140 3.810 12.700 4.050 ;
        RECT  14.790 1.630 15.030 4.350 ;
        RECT  15.850 1.860 16.840 2.100 ;
        RECT  16.600 2.440 17.230 2.680 ;
        RECT  16.600 1.860 16.840 3.530 ;
        RECT  15.780 3.290 16.840 3.530 ;
        RECT  5.390 1.130 18.230 1.370 ;
        RECT  17.710 0.980 18.230 1.400 ;
        RECT  11.820 1.130 12.060 2.900 ;
        RECT  17.990 0.980 18.230 3.470 ;
        RECT  11.960 2.600 12.200 3.570 ;
        RECT  5.390 1.130 5.630 3.650 ;
        RECT  5.170 3.250 5.630 3.650 ;
        RECT  17.180 1.780 17.710 2.180 ;
        RECT  17.080 3.290 17.710 3.530 ;
        RECT  17.470 1.780 17.710 4.020 ;
        RECT  17.470 3.780 18.490 4.020 ;
        RECT  19.230 1.450 19.540 3.470 ;
        RECT  19.230 3.070 19.710 3.470 ;
        RECT  18.560 1.450 18.800 2.700 ;
        RECT  19.950 2.620 20.860 2.860 ;
        RECT  18.730 2.400 18.970 3.950 ;
        RECT  19.950 2.620 20.190 3.950 ;
        RECT  18.730 3.710 20.190 3.950 ;
        RECT  20.790 1.450 21.030 2.300 ;
        RECT  19.780 2.060 21.390 2.300 ;
        RECT  21.150 2.060 21.390 3.390 ;
        RECT  20.820 3.150 21.390 3.390 ;
        RECT  22.280 1.480 22.520 3.950 ;
        RECT  22.280 3.160 22.760 3.950 ;
        RECT  20.430 3.710 22.760 3.950 ;
        RECT  15.270 3.420 15.510 4.370 ;
        RECT  18.660 4.190 20.670 4.430 ;
        RECT  15.270 4.130 17.250 4.370 ;
        RECT  20.430 3.710 20.670 4.430 ;
        RECT  17.010 4.300 18.900 4.540 ;
        RECT  21.520 1.000 23.000 1.240 ;
        RECT  21.520 1.000 21.930 1.850 ;
        RECT  22.760 1.000 23.000 2.380 ;
        RECT  22.760 2.140 23.970 2.380 ;
        RECT  21.690 1.000 21.930 3.470 ;
        RECT  23.860 1.610 24.450 1.850 ;
        RECT  24.210 1.610 24.450 2.860 ;
        RECT  24.210 2.610 25.150 2.860 ;
        RECT  22.760 2.620 25.150 2.860 ;
        RECT  23.900 2.620 24.140 3.470 ;
    END
END senrq1

MACRO senrb4
    CLASS CORE ;
    FOREIGN senrb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 2.020 8.900 2.460 ;
        RECT  8.350 2.200 8.750 2.600 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 4.980 2.460 ;
        RECT  4.140 2.040 4.980 2.440 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.880 2.510 6.320 2.910 ;
        RECT  5.880 1.970 6.120 2.910 ;
        RECT  5.220 1.970 6.120 2.210 ;
        RECT  5.220 1.540 5.460 2.210 ;
        RECT  4.020 1.540 5.460 1.780 ;
        RECT  3.060 1.460 4.260 1.700 ;
        RECT  3.060 1.460 3.300 2.460 ;
        RECT  2.760 2.220 3.160 2.810 ;
        RECT  2.860 2.020 3.300 2.460 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.218  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  21.600 1.100 22.020 1.520 ;
        RECT  19.540 3.930 21.810 4.330 ;
        RECT  21.340 1.230 21.810 4.330 ;
        RECT  20.460 1.230 22.020 1.470 ;
        RECT  20.080 1.200 20.620 1.440 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.039  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.380 1.200 19.000 1.440 ;
        RECT  16.890 2.990 18.630 3.390 ;
        RECT  17.380 1.220 18.570 1.460 ;
        RECT  17.980 1.220 18.420 3.390 ;
        RECT  17.120 0.980 17.620 1.300 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.449  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.710 0.540 3.110 ;
        RECT  0.120 2.020 0.500 2.880 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.387  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.020 7.780 2.460 ;
        RECT  7.170 2.030 7.780 2.430 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 22.400 5.600 ;
        RECT  21.590 4.620 21.990 5.600 ;
        RECT  20.280 4.620 20.680 5.600 ;
        RECT  18.970 4.620 19.370 5.600 ;
        RECT  17.630 4.550 18.030 5.600 ;
        RECT  16.320 4.110 16.720 5.600 ;
        RECT  14.920 4.620 15.320 5.600 ;
        RECT  12.280 4.710 12.600 5.600 ;
        RECT  8.920 4.710 9.320 5.600 ;
        RECT  6.180 4.620 6.580 5.600 ;
        RECT  2.810 4.370 3.320 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 22.400 0.740 ;
        RECT  20.820 0.000 21.220 0.990 ;
        RECT  19.340 0.000 19.740 0.980 ;
        RECT  17.860 0.000 18.260 0.980 ;
        RECT  15.720 0.000 16.040 0.980 ;
        RECT  12.590 0.000 12.990 0.890 ;
        RECT  8.890 0.000 9.290 0.890 ;
        RECT  6.280 0.000 6.680 1.200 ;
        RECT  2.410 0.000 2.830 0.930 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.420 0.980 1.660 ;
        RECT  0.740 1.420 0.980 2.240 ;
        RECT  0.740 2.000 1.260 2.240 ;
        RECT  1.020 2.000 1.260 3.690 ;
        RECT  0.150 3.450 1.260 3.690 ;
        RECT  1.220 0.980 1.940 1.220 ;
        RECT  1.220 0.980 1.460 1.710 ;
        RECT  1.220 1.470 1.740 1.710 ;
        RECT  1.500 1.470 1.740 2.490 ;
        RECT  1.500 2.250 2.030 2.490 ;
        RECT  1.790 2.250 2.030 2.980 ;
        RECT  1.570 2.740 1.810 3.680 ;
        RECT  2.060 1.590 2.520 1.990 ;
        RECT  3.540 2.180 3.780 3.360 ;
        RECT  2.280 3.120 3.780 3.360 ;
        RECT  2.280 1.590 2.520 3.620 ;
        RECT  2.200 3.380 2.440 4.480 ;
        RECT  8.280 1.540 9.380 1.780 ;
        RECT  9.140 2.100 9.620 2.500 ;
        RECT  9.140 1.540 9.380 2.670 ;
        RECT  9.120 2.560 9.360 3.210 ;
        RECT  8.230 2.970 9.360 3.210 ;
        RECT  9.720 1.210 9.960 1.880 ;
        RECT  9.720 1.640 10.220 1.880 ;
        RECT  9.980 1.640 10.220 2.490 ;
        RECT  9.860 2.280 10.100 2.990 ;
        RECT  9.610 2.750 10.100 2.990 ;
        RECT  9.610 2.750 9.850 3.310 ;
        RECT  4.330 0.980 5.390 1.220 ;
        RECT  5.170 1.060 5.940 1.300 ;
        RECT  10.340 0.980 10.740 1.380 ;
        RECT  6.920 1.170 7.880 1.410 ;
        RECT  5.700 1.060 5.940 1.730 ;
        RECT  6.920 1.170 7.160 1.730 ;
        RECT  5.700 1.490 7.160 1.730 ;
        RECT  10.500 0.980 10.740 2.590 ;
        RECT  10.500 0.980 10.700 2.930 ;
        RECT  6.560 1.490 6.800 3.700 ;
        RECT  10.460 2.450 10.580 4.050 ;
        RECT  10.340 2.710 10.580 4.050 ;
        RECT  5.020 3.460 7.990 3.700 ;
        RECT  4.540 3.560 5.260 3.800 ;
        RECT  7.750 3.560 8.920 3.800 ;
        RECT  8.680 3.740 10.580 3.980 ;
        RECT  10.130 3.650 10.580 4.050 ;
        RECT  11.660 1.650 12.220 1.890 ;
        RECT  11.660 1.650 11.900 2.150 ;
        RECT  11.460 1.910 11.700 3.730 ;
        RECT  11.550 3.490 11.790 4.050 ;
        RECT  10.980 1.130 12.980 1.410 ;
        RECT  10.980 1.130 11.480 1.480 ;
        RECT  10.980 1.130 11.400 1.560 ;
        RECT  12.740 1.130 12.980 2.810 ;
        RECT  10.980 1.130 11.220 3.460 ;
        RECT  10.820 3.140 11.220 3.460 ;
        RECT  13.310 0.980 13.760 1.300 ;
        RECT  11.940 2.560 12.180 3.130 ;
        RECT  13.310 0.980 13.550 3.220 ;
        RECT  12.150 2.890 12.390 3.990 ;
        RECT  13.140 2.990 13.380 3.990 ;
        RECT  12.150 3.750 13.380 3.990 ;
        RECT  13.830 1.540 14.070 2.220 ;
        RECT  13.870 1.980 14.110 3.060 ;
        RECT  14.950 1.600 15.190 2.230 ;
        RECT  5.240 2.460 5.640 2.860 ;
        RECT  4.030 2.720 5.450 2.960 ;
        RECT  4.030 2.720 4.520 3.120 ;
        RECT  14.910 1.940 15.150 4.170 ;
        RECT  4.030 2.720 4.270 4.280 ;
        RECT  14.280 3.930 15.150 4.170 ;
        RECT  4.030 4.040 8.440 4.280 ;
        RECT  8.200 4.230 9.800 4.470 ;
        RECT  11.950 4.230 13.200 4.470 ;
        RECT  9.560 4.290 12.110 4.530 ;
        RECT  14.280 3.930 14.680 4.620 ;
        RECT  12.960 4.380 14.680 4.620 ;
        RECT  14.100 1.170 15.550 1.300 ;
        RECT  14.100 1.060 14.650 1.300 ;
        RECT  14.430 1.120 15.500 1.360 ;
        RECT  15.350 1.220 16.200 1.420 ;
        RECT  15.400 1.220 16.200 1.460 ;
        RECT  15.960 1.220 16.200 2.270 ;
        RECT  15.960 1.870 16.510 2.270 ;
        RECT  14.430 1.120 14.670 3.690 ;
        RECT  13.620 3.450 14.670 3.690 ;
        RECT  13.620 3.450 13.860 4.070 ;
        RECT  16.460 1.450 16.930 1.630 ;
        RECT  16.460 0.980 16.700 1.630 ;
        RECT  16.680 1.390 16.850 1.700 ;
        RECT  15.480 1.700 15.720 2.750 ;
        RECT  16.750 1.530 16.990 2.750 ;
        RECT  15.480 2.510 16.990 2.750 ;
        RECT  19.000 2.350 20.770 2.750 ;
        RECT  15.700 2.510 15.940 3.870 ;
        RECT  19.000 2.350 19.240 3.870 ;
        RECT  15.700 3.630 19.240 3.870 ;
    END
END senrb4

MACRO senrb2
    CLASS CORE ;
    FOREIGN senrb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 2.020 8.900 2.460 ;
        RECT  8.350 2.200 8.750 2.600 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 4.980 2.460 ;
        RECT  4.140 2.040 4.980 2.440 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.880 2.510 6.320 2.910 ;
        RECT  5.880 1.970 6.120 2.910 ;
        RECT  5.220 1.970 6.120 2.210 ;
        RECT  5.220 1.540 5.460 2.210 ;
        RECT  4.020 1.540 5.460 1.780 ;
        RECT  3.060 1.460 4.260 1.700 ;
        RECT  3.060 1.460 3.300 2.460 ;
        RECT  2.760 2.220 3.160 2.810 ;
        RECT  2.860 2.020 3.300 2.460 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.920  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.470 3.930 19.480 4.330 ;
        RECT  19.100 1.880 19.480 4.330 ;
        RECT  19.050 1.500 19.450 2.020 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.796  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.300 1.980 17.860 2.490 ;
        RECT  16.890 2.930 17.700 3.260 ;
        RECT  17.300 1.680 17.700 3.260 ;
        RECT  17.110 1.680 17.700 2.080 ;
        RECT  16.890 2.930 17.290 3.500 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.449  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.710 0.540 3.110 ;
        RECT  0.120 2.020 0.500 2.880 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.387  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.020 7.780 2.460 ;
        RECT  7.170 2.030 7.780 2.430 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.600 5.600 ;
        RECT  19.040 4.620 19.440 5.600 ;
        RECT  17.630 4.620 18.030 5.600 ;
        RECT  16.320 4.620 16.730 5.600 ;
        RECT  14.920 4.620 15.320 5.600 ;
        RECT  12.280 4.710 12.600 5.600 ;
        RECT  8.920 4.710 9.320 5.600 ;
        RECT  6.180 4.620 6.580 5.600 ;
        RECT  2.810 4.370 3.320 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.600 0.740 ;
        RECT  18.310 0.000 18.710 0.980 ;
        RECT  15.720 0.000 16.040 0.980 ;
        RECT  12.590 0.000 12.990 0.890 ;
        RECT  8.890 0.000 9.290 0.890 ;
        RECT  6.280 0.000 6.680 1.200 ;
        RECT  2.410 0.000 2.830 0.930 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.420 0.980 1.660 ;
        RECT  0.740 1.420 0.980 2.240 ;
        RECT  0.740 2.000 1.260 2.240 ;
        RECT  1.020 2.000 1.260 3.690 ;
        RECT  0.150 3.450 1.260 3.690 ;
        RECT  1.220 0.980 1.940 1.220 ;
        RECT  1.220 0.980 1.460 1.710 ;
        RECT  1.220 1.470 1.740 1.710 ;
        RECT  1.500 1.470 1.740 2.490 ;
        RECT  1.500 2.250 2.030 2.490 ;
        RECT  1.790 2.250 2.030 2.980 ;
        RECT  1.570 2.740 1.810 3.680 ;
        RECT  2.060 1.590 2.520 1.990 ;
        RECT  3.540 2.180 3.780 3.360 ;
        RECT  2.280 3.120 3.780 3.360 ;
        RECT  2.280 1.590 2.520 3.620 ;
        RECT  2.200 3.380 2.440 4.480 ;
        RECT  8.280 1.540 9.380 1.780 ;
        RECT  9.140 2.100 9.620 2.500 ;
        RECT  9.140 1.540 9.380 2.670 ;
        RECT  9.120 2.560 9.360 3.210 ;
        RECT  8.230 2.970 9.360 3.210 ;
        RECT  9.720 1.210 9.960 1.880 ;
        RECT  9.720 1.640 10.220 1.880 ;
        RECT  9.980 1.640 10.220 2.490 ;
        RECT  9.860 2.280 10.100 2.990 ;
        RECT  9.610 2.750 10.100 2.990 ;
        RECT  9.610 2.750 9.850 3.310 ;
        RECT  4.330 0.980 5.390 1.220 ;
        RECT  5.170 1.060 5.940 1.300 ;
        RECT  10.340 0.980 10.740 1.380 ;
        RECT  6.920 1.170 7.880 1.410 ;
        RECT  5.700 1.060 5.940 1.730 ;
        RECT  6.920 1.170 7.160 1.730 ;
        RECT  5.700 1.490 7.160 1.730 ;
        RECT  10.500 0.980 10.740 2.590 ;
        RECT  10.500 0.980 10.700 2.930 ;
        RECT  6.560 1.490 6.800 3.700 ;
        RECT  10.460 2.450 10.580 4.050 ;
        RECT  10.340 2.710 10.580 4.050 ;
        RECT  5.020 3.460 7.990 3.700 ;
        RECT  4.540 3.560 5.260 3.800 ;
        RECT  7.750 3.560 8.920 3.800 ;
        RECT  8.680 3.740 10.580 3.980 ;
        RECT  10.130 3.650 10.580 4.050 ;
        RECT  11.660 1.650 12.220 1.890 ;
        RECT  11.660 1.650 11.900 2.150 ;
        RECT  11.460 1.910 11.700 3.730 ;
        RECT  11.550 3.490 11.790 4.050 ;
        RECT  10.980 1.130 12.980 1.410 ;
        RECT  10.980 1.130 11.480 1.480 ;
        RECT  10.980 1.130 11.400 1.560 ;
        RECT  12.740 1.130 12.980 2.810 ;
        RECT  10.980 1.130 11.220 3.460 ;
        RECT  10.820 3.140 11.220 3.460 ;
        RECT  13.310 0.980 13.760 1.300 ;
        RECT  11.940 2.560 12.180 3.130 ;
        RECT  13.310 0.980 13.550 3.220 ;
        RECT  12.150 2.890 12.390 3.990 ;
        RECT  13.140 2.990 13.380 3.990 ;
        RECT  12.150 3.750 13.380 3.990 ;
        RECT  13.830 1.540 14.070 2.220 ;
        RECT  13.870 1.980 14.110 3.060 ;
        RECT  14.950 1.600 15.190 2.230 ;
        RECT  5.240 2.460 5.640 2.860 ;
        RECT  4.030 2.720 5.450 2.960 ;
        RECT  4.030 2.720 4.520 3.120 ;
        RECT  14.910 1.940 15.150 4.170 ;
        RECT  4.030 2.720 4.270 4.280 ;
        RECT  14.280 3.930 15.150 4.170 ;
        RECT  4.030 4.040 8.440 4.280 ;
        RECT  8.200 4.230 9.800 4.470 ;
        RECT  11.950 4.230 13.200 4.470 ;
        RECT  9.560 4.290 12.110 4.530 ;
        RECT  14.280 3.930 14.680 4.620 ;
        RECT  12.960 4.380 14.680 4.620 ;
        RECT  14.100 1.170 15.550 1.300 ;
        RECT  14.100 1.060 14.650 1.300 ;
        RECT  14.430 1.120 15.500 1.360 ;
        RECT  15.350 1.220 16.200 1.420 ;
        RECT  15.400 1.220 16.200 1.460 ;
        RECT  15.960 1.220 16.200 2.690 ;
        RECT  15.960 2.290 16.980 2.690 ;
        RECT  14.430 1.120 14.670 3.690 ;
        RECT  13.620 3.450 14.670 3.690 ;
        RECT  13.620 3.450 13.860 4.070 ;
        RECT  16.490 1.080 18.080 1.320 ;
        RECT  17.840 1.240 18.710 1.480 ;
        RECT  16.490 1.080 16.730 1.800 ;
        RECT  15.480 1.700 15.720 2.750 ;
        RECT  15.440 2.510 15.680 3.350 ;
        RECT  15.440 3.110 16.200 3.350 ;
        RECT  18.470 1.240 18.710 3.640 ;
        RECT  17.900 3.400 18.710 3.640 ;
        RECT  15.960 3.110 16.200 4.220 ;
        RECT  17.900 3.400 18.140 4.220 ;
        RECT  15.960 3.980 18.140 4.220 ;
    END
END senrb2

MACRO senrb1
    CLASS CORE ;
    FOREIGN senrb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 2.020 8.900 2.460 ;
        RECT  8.350 2.200 8.750 2.600 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 4.980 2.460 ;
        RECT  4.140 2.040 4.980 2.440 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.880 2.510 6.320 2.910 ;
        RECT  5.880 1.970 6.120 2.910 ;
        RECT  5.220 1.970 6.120 2.210 ;
        RECT  5.220 1.540 5.460 2.210 ;
        RECT  4.020 1.540 5.460 1.780 ;
        RECT  3.060 1.460 4.260 1.700 ;
        RECT  3.060 1.460 3.300 2.460 ;
        RECT  2.760 2.220 3.160 2.810 ;
        RECT  2.860 2.020 3.300 2.460 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.170  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.420 1.980 17.860 2.490 ;
        RECT  17.310 2.480 17.700 2.720 ;
        RECT  17.080 1.810 17.660 2.050 ;
        RECT  16.970 2.930 17.550 3.170 ;
        RECT  17.310 2.480 17.550 3.170 ;
        RECT  16.510 3.730 17.210 3.980 ;
        RECT  16.970 2.930 17.210 3.980 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.345  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.980 2.960 18.760 3.200 ;
        RECT  18.520 1.040 18.760 3.200 ;
        RECT  17.850 3.460 18.420 3.860 ;
        RECT  17.980 2.960 18.420 3.860 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.449  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.710 0.540 3.110 ;
        RECT  0.120 2.020 0.500 2.880 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.387  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.020 7.780 2.460 ;
        RECT  7.170 2.030 7.780 2.430 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.040 5.600 ;
        RECT  17.220 4.620 17.620 5.600 ;
        RECT  15.000 4.620 15.400 5.600 ;
        RECT  12.290 4.710 12.690 5.600 ;
        RECT  8.920 4.710 9.320 5.600 ;
        RECT  6.180 4.620 6.580 5.600 ;
        RECT  2.810 4.370 3.320 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.040 0.740 ;
        RECT  17.460 0.000 17.860 0.980 ;
        RECT  15.720 0.000 15.960 0.980 ;
        RECT  12.590 0.000 12.990 0.890 ;
        RECT  9.050 0.000 9.450 0.890 ;
        RECT  6.280 0.000 6.680 1.200 ;
        RECT  2.410 0.000 2.830 0.930 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.420 0.980 1.660 ;
        RECT  0.740 1.420 0.980 2.240 ;
        RECT  0.740 2.000 1.260 2.240 ;
        RECT  1.020 2.000 1.260 3.690 ;
        RECT  0.150 3.450 1.260 3.690 ;
        RECT  1.220 0.980 1.940 1.220 ;
        RECT  1.220 0.980 1.460 1.710 ;
        RECT  1.220 1.470 1.740 1.710 ;
        RECT  1.500 1.470 1.740 2.490 ;
        RECT  1.500 2.250 2.030 2.490 ;
        RECT  1.790 2.250 2.030 2.980 ;
        RECT  1.570 2.740 1.810 3.680 ;
        RECT  2.060 1.590 2.520 1.990 ;
        RECT  3.540 2.180 3.780 3.360 ;
        RECT  2.280 3.120 3.780 3.360 ;
        RECT  2.280 1.590 2.520 3.620 ;
        RECT  2.200 3.380 2.440 4.480 ;
        RECT  8.280 1.540 9.380 1.780 ;
        RECT  9.140 1.540 9.380 2.670 ;
        RECT  9.140 2.180 9.620 2.600 ;
        RECT  9.120 2.560 9.440 2.670 ;
        RECT  9.120 2.560 9.360 3.210 ;
        RECT  8.230 2.970 9.360 3.210 ;
        RECT  9.720 1.300 9.960 1.940 ;
        RECT  9.720 1.700 10.220 1.940 ;
        RECT  9.980 1.700 10.220 3.180 ;
        RECT  9.610 2.940 10.220 3.180 ;
        RECT  9.610 2.940 9.850 3.510 ;
        RECT  4.330 0.980 5.390 1.220 ;
        RECT  5.170 1.060 5.940 1.300 ;
        RECT  10.340 0.980 10.740 1.380 ;
        RECT  6.920 1.170 7.880 1.410 ;
        RECT  5.700 1.060 5.940 1.730 ;
        RECT  6.920 1.170 7.160 1.730 ;
        RECT  5.700 1.490 7.160 1.730 ;
        RECT  6.560 1.490 6.800 3.700 ;
        RECT  5.020 3.460 7.990 3.700 ;
        RECT  4.540 3.560 5.260 3.800 ;
        RECT  7.750 3.560 8.920 3.800 ;
        RECT  8.680 3.750 10.740 3.990 ;
        RECT  10.500 0.980 10.740 4.080 ;
        RECT  10.300 3.750 10.740 4.080 ;
        RECT  11.660 1.650 12.220 1.890 ;
        RECT  11.660 1.650 11.900 2.150 ;
        RECT  11.540 1.910 11.780 3.570 ;
        RECT  11.670 3.330 11.910 3.970 ;
        RECT  10.980 1.130 13.070 1.410 ;
        RECT  10.980 1.130 11.480 1.480 ;
        RECT  10.980 1.130 11.400 1.560 ;
        RECT  12.830 1.130 13.070 2.570 ;
        RECT  10.980 1.130 11.220 3.400 ;
        RECT  13.310 0.980 13.790 1.300 ;
        RECT  13.310 0.980 13.550 3.080 ;
        RECT  12.020 2.470 12.260 3.090 ;
        RECT  12.150 2.850 12.390 3.640 ;
        RECT  13.260 2.820 13.500 3.640 ;
        RECT  12.150 3.400 13.500 3.640 ;
        RECT  12.970 3.400 13.210 3.970 ;
        RECT  13.830 1.540 14.070 2.220 ;
        RECT  13.950 1.980 14.190 3.060 ;
        RECT  14.950 1.620 15.190 2.230 ;
        RECT  5.240 2.460 5.640 2.860 ;
        RECT  4.030 2.720 5.450 2.960 ;
        RECT  4.030 2.720 4.520 3.120 ;
        RECT  14.910 1.940 15.150 4.020 ;
        RECT  14.480 3.780 15.150 4.020 ;
        RECT  4.030 2.720 4.270 4.280 ;
        RECT  4.030 4.040 8.440 4.280 ;
        RECT  8.200 4.230 10.060 4.470 ;
        RECT  10.980 4.230 13.200 4.470 ;
        RECT  9.820 4.320 11.220 4.560 ;
        RECT  14.480 3.780 14.720 4.620 ;
        RECT  12.960 4.380 14.720 4.620 ;
        RECT  14.100 1.060 14.650 1.300 ;
        RECT  14.430 1.140 15.530 1.380 ;
        RECT  15.350 1.220 16.250 1.430 ;
        RECT  15.400 1.220 16.250 1.460 ;
        RECT  16.010 1.220 16.250 2.770 ;
        RECT  14.430 1.140 14.670 3.540 ;
        RECT  13.740 3.300 14.670 3.540 ;
        RECT  13.740 3.300 13.980 3.970 ;
        RECT  16.490 2.290 17.060 2.690 ;
        RECT  15.490 1.700 15.730 2.710 ;
        RECT  15.420 2.470 15.660 3.360 ;
        RECT  16.490 0.990 16.730 3.360 ;
        RECT  15.420 3.120 16.730 3.360 ;
    END
END senrb1

MACRO secrq4
    CLASS CORE ;
    FOREIGN secrq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.910 2.400 17.390 2.800 ;
        RECT  16.910 2.400 17.220 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.690 2.020 11.930 2.770 ;
        RECT  11.260 2.020 11.930 2.460 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.530 3.140 4.980 3.580 ;
        RECT  4.530 2.600 4.770 3.580 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.458  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.400 2.020 7.360 2.460 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.261  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.390 1.740 21.130 1.980 ;
        RECT  20.070 2.560 20.670 3.020 ;
        RECT  19.990 3.830 20.400 4.260 ;
        RECT  20.070 1.740 20.400 4.260 ;
        RECT  18.760 3.970 20.400 4.210 ;
        RECT  18.760 3.630 19.000 4.210 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.533  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.420 0.570 2.820 ;
        RECT  0.120 2.020 0.500 2.820 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.362  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.620 2.000 4.390 2.240 ;
        RECT  3.620 1.460 3.860 2.240 ;
        RECT  3.420 1.460 3.860 1.900 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 21.280 5.600 ;
        RECT  20.730 4.550 21.130 5.600 ;
        RECT  19.420 4.550 19.820 5.600 ;
        RECT  18.110 4.370 18.510 5.600 ;
        RECT  16.760 4.520 17.160 5.600 ;
        RECT  14.190 4.710 14.590 5.600 ;
        RECT  11.760 4.710 12.160 5.600 ;
        RECT  10.420 4.710 10.820 5.600 ;
        RECT  6.300 4.620 6.700 5.600 ;
        RECT  2.800 4.620 3.200 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 21.280 0.740 ;
        RECT  19.970 0.000 20.370 1.180 ;
        RECT  16.850 0.000 17.250 1.680 ;
        RECT  13.240 0.000 13.640 1.280 ;
        RECT  11.210 0.000 11.450 1.280 ;
        RECT  9.100 0.000 9.500 0.820 ;
        RECT  6.460 0.000 6.700 1.230 ;
        RECT  2.180 0.000 2.580 1.020 ;
        RECT  0.890 0.000 1.290 1.020 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 0.980 0.470 1.580 ;
        RECT  0.230 1.340 1.160 1.580 ;
        RECT  0.920 1.340 1.160 2.630 ;
        RECT  0.810 2.390 1.050 3.300 ;
        RECT  2.800 2.980 3.560 3.220 ;
        RECT  0.230 3.060 1.050 3.300 ;
        RECT  0.230 3.060 0.470 4.370 ;
        RECT  2.800 2.980 3.040 4.370 ;
        RECT  0.230 4.130 3.040 4.370 ;
        RECT  2.930 0.980 4.470 1.220 ;
        RECT  2.930 0.980 3.170 1.500 ;
        RECT  1.590 1.260 3.170 1.500 ;
        RECT  4.230 0.980 4.470 1.760 ;
        RECT  4.230 1.520 5.260 1.760 ;
        RECT  1.590 1.260 1.830 2.310 ;
        RECT  5.020 1.520 5.260 2.900 ;
        RECT  1.400 2.070 1.640 3.300 ;
        RECT  5.220 2.660 5.460 3.420 ;
        RECT  5.220 3.180 6.610 3.420 ;
        RECT  1.330 3.060 1.570 3.890 ;
        RECT  1.330 3.650 1.930 3.890 ;
        RECT  5.660 1.980 6.160 2.380 ;
        RECT  2.290 1.740 2.530 2.730 ;
        RECT  5.920 1.980 6.160 2.940 ;
        RECT  2.290 2.490 4.040 2.730 ;
        RECT  5.920 2.700 7.430 2.940 ;
        RECT  2.310 2.490 2.550 3.850 ;
        RECT  3.800 2.490 4.040 4.140 ;
        RECT  5.340 3.660 7.430 3.900 ;
        RECT  7.190 2.700 7.430 3.900 ;
        RECT  3.800 3.900 5.580 4.140 ;
        RECT  7.670 0.980 8.720 1.220 ;
        RECT  4.710 1.040 6.220 1.280 ;
        RECT  5.980 1.040 6.220 1.710 ;
        RECT  6.940 1.410 7.910 1.650 ;
        RECT  5.980 1.470 7.180 1.710 ;
        RECT  7.670 0.980 7.910 4.460 ;
        RECT  5.820 4.140 7.200 4.380 ;
        RECT  6.960 4.220 8.460 4.460 ;
        RECT  4.300 4.380 6.060 4.620 ;
        RECT  9.970 1.840 10.210 2.660 ;
        RECT  9.660 2.420 10.210 2.660 ;
        RECT  9.660 2.420 9.900 3.420 ;
        RECT  9.540 3.180 9.780 3.900 ;
        RECT  9.540 3.660 11.470 3.900 ;
        RECT  12.170 1.800 12.410 2.620 ;
        RECT  12.170 2.380 12.920 2.620 ;
        RECT  12.630 2.380 12.920 2.940 ;
        RECT  12.680 2.380 12.920 3.500 ;
        RECT  12.340 3.260 12.920 3.500 ;
        RECT  8.630 1.940 9.490 2.180 ;
        RECT  8.630 1.940 8.870 2.660 ;
        RECT  8.630 2.420 9.280 2.660 ;
        RECT  9.040 2.420 9.280 4.470 ;
        RECT  9.040 4.230 12.540 4.470 ;
        RECT  13.870 4.230 14.440 4.470 ;
        RECT  14.200 2.630 14.440 4.470 ;
        RECT  12.320 4.290 14.030 4.530 ;
        RECT  13.640 2.140 14.830 2.380 ;
        RECT  14.360 1.790 14.600 2.380 ;
        RECT  14.580 2.220 14.940 2.430 ;
        RECT  10.140 2.900 11.450 3.140 ;
        RECT  11.210 3.020 11.950 3.260 ;
        RECT  11.710 3.020 11.950 3.990 ;
        RECT  11.710 3.740 12.960 3.990 ;
        RECT  13.550 3.760 13.880 3.990 ;
        RECT  14.700 2.220 14.940 3.810 ;
        RECT  13.640 2.140 13.880 3.990 ;
        RECT  12.710 3.810 13.710 4.050 ;
        RECT  11.690 0.990 12.980 1.230 ;
        RECT  8.960 1.060 10.770 1.300 ;
        RECT  14.850 1.110 15.900 1.350 ;
        RECT  13.880 1.120 14.930 1.360 ;
        RECT  10.530 1.060 10.770 1.760 ;
        RECT  12.740 0.990 12.980 2.020 ;
        RECT  8.960 1.060 9.200 1.700 ;
        RECT  8.150 1.460 9.200 1.700 ;
        RECT  11.690 0.990 11.930 1.760 ;
        RECT  10.530 1.520 11.930 1.760 ;
        RECT  13.880 1.120 14.120 1.860 ;
        RECT  12.740 1.620 14.120 1.860 ;
        RECT  12.740 1.620 13.400 2.020 ;
        RECT  15.660 1.110 15.900 3.270 ;
        RECT  8.150 1.460 8.390 3.140 ;
        RECT  8.150 2.900 8.700 3.140 ;
        RECT  15.660 2.870 16.060 3.270 ;
        RECT  13.160 1.620 13.400 3.570 ;
        RECT  15.020 1.590 15.420 1.990 ;
        RECT  17.750 2.600 17.990 3.500 ;
        RECT  16.830 3.260 17.990 3.500 ;
        RECT  15.180 1.590 15.420 4.390 ;
        RECT  15.790 4.040 17.070 4.280 ;
        RECT  16.830 3.260 17.070 4.280 ;
        RECT  15.180 4.150 16.030 4.390 ;
        RECT  17.490 0.980 19.000 1.220 ;
        RECT  17.490 0.980 17.730 2.160 ;
        RECT  16.140 1.920 17.730 2.160 ;
        RECT  16.140 1.580 16.380 2.230 ;
        RECT  16.350 1.920 16.590 3.780 ;
        RECT  16.020 3.540 16.590 3.780 ;
        RECT  18.050 1.620 18.910 1.860 ;
        RECT  18.670 2.390 19.620 2.790 ;
        RECT  18.670 1.620 18.910 3.390 ;
        RECT  18.280 3.150 18.910 3.390 ;
        RECT  18.280 3.150 18.520 3.980 ;
        RECT  17.360 3.740 18.520 3.980 ;
    END
END secrq4

MACRO secrq2
    CLASS CORE ;
    FOREIGN secrq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.440 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.419  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  24.720 2.400 25.130 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.405  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.720 2.510 16.330 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.940 2.250 13.380 3.020 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.397  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.700 2.580 7.310 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.177  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  26.240 3.110 26.740 3.510 ;
        RECT  26.460 1.480 26.740 3.510 ;
        RECT  26.300 1.480 26.740 1.880 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.020 0.980 2.900 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.280 1.640 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 27.440 5.600 ;
        RECT  26.880 4.190 27.120 5.600 ;
        RECT  25.540 4.190 25.780 5.600 ;
        RECT  24.240 4.190 24.480 5.600 ;
        RECT  20.080 4.580 20.480 5.600 ;
        RECT  16.280 4.710 16.680 5.600 ;
        RECT  14.640 4.710 15.040 5.600 ;
        RECT  13.390 4.710 13.790 5.600 ;
        RECT  9.670 4.480 10.070 5.600 ;
        RECT  8.200 3.770 8.440 5.600 ;
        RECT  6.900 3.770 7.140 5.600 ;
        RECT  6.000 3.850 6.240 5.600 ;
        RECT  3.930 4.090 4.170 5.600 ;
        RECT  1.660 4.460 2.060 5.600 ;
        RECT  0.970 3.290 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 27.440 0.740 ;
        RECT  26.970 0.000 27.210 1.210 ;
        RECT  25.640 0.000 25.880 1.300 ;
        RECT  20.470 0.000 20.710 1.980 ;
        RECT  16.460 0.000 16.860 0.890 ;
        RECT  15.050 0.000 15.450 0.890 ;
        RECT  13.070 0.000 13.470 0.890 ;
        RECT  10.170 0.000 10.570 0.890 ;
        RECT  8.130 0.000 8.530 0.890 ;
        RECT  6.180 0.000 6.600 0.890 ;
        RECT  4.190 0.000 4.430 1.470 ;
        RECT  1.660 0.000 2.060 1.140 ;
        RECT  0.760 0.000 1.180 1.180 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 1.520 0.470 1.920 ;
        RECT  0.220 1.520 0.460 4.620 ;
        RECT  0.220 3.290 0.470 4.620 ;
        RECT  1.570 1.530 2.120 1.850 ;
        RECT  1.880 2.270 2.990 2.510 ;
        RECT  1.880 1.530 2.120 3.650 ;
        RECT  1.630 3.330 2.120 3.650 ;
        RECT  2.430 0.980 2.990 1.300 ;
        RECT  2.670 0.980 2.990 1.910 ;
        RECT  2.670 1.630 3.470 1.910 ;
        RECT  3.230 1.630 3.470 2.990 ;
        RECT  2.480 2.750 3.470 2.990 ;
        RECT  2.480 2.750 2.720 4.620 ;
        RECT  2.430 4.220 2.830 4.620 ;
        RECT  3.230 1.150 3.950 1.390 ;
        RECT  3.710 2.800 4.450 3.040 ;
        RECT  3.710 1.150 3.950 3.610 ;
        RECT  2.960 3.370 3.950 3.610 ;
        RECT  2.960 3.370 3.280 3.770 ;
        RECT  4.570 1.830 4.930 2.150 ;
        RECT  4.690 1.830 4.930 3.750 ;
        RECT  4.430 3.430 4.930 3.750 ;
        RECT  6.000 1.610 6.580 1.850 ;
        RECT  6.000 1.610 6.240 3.510 ;
        RECT  9.440 1.610 9.680 2.500 ;
        RECT  9.160 2.260 10.280 2.500 ;
        RECT  9.160 2.260 9.400 3.740 ;
        RECT  10.170 1.690 10.760 1.930 ;
        RECT  10.520 1.690 10.760 3.740 ;
        RECT  10.520 2.510 11.050 2.910 ;
        RECT  10.520 2.510 10.840 3.740 ;
        RECT  10.440 3.340 10.840 3.740 ;
        RECT  12.460 1.610 12.880 1.930 ;
        RECT  12.460 1.610 12.700 3.510 ;
        RECT  12.460 3.270 13.020 3.510 ;
        RECT  6.900 1.620 7.860 1.860 ;
        RECT  7.620 1.620 7.860 3.510 ;
        RECT  7.540 3.110 7.940 3.510 ;
        RECT  7.540 3.270 8.920 3.510 ;
        RECT  8.680 3.270 8.920 4.240 ;
        RECT  8.680 4.000 10.600 4.240 ;
        RECT  10.360 4.000 10.600 4.530 ;
        RECT  12.900 4.230 14.140 4.470 ;
        RECT  10.360 4.290 13.140 4.530 ;
        RECT  13.930 1.610 14.170 2.540 ;
        RECT  13.930 2.140 14.530 2.540 ;
        RECT  14.070 2.140 14.310 3.510 ;
        RECT  11.000 1.610 11.540 1.930 ;
        RECT  14.790 1.710 15.450 1.950 ;
        RECT  11.300 1.610 11.540 4.050 ;
        RECT  11.140 3.250 11.540 4.050 ;
        RECT  12.400 3.750 15.030 3.990 ;
        RECT  11.140 3.810 12.700 4.050 ;
        RECT  14.790 1.710 15.030 4.350 ;
        RECT  15.850 1.910 16.810 2.150 ;
        RECT  16.570 2.760 17.180 3.000 ;
        RECT  16.570 1.910 16.810 3.530 ;
        RECT  15.750 3.290 16.810 3.530 ;
        RECT  17.150 1.830 17.660 2.230 ;
        RECT  17.050 3.290 17.660 3.530 ;
        RECT  17.420 1.830 17.660 4.140 ;
        RECT  17.420 3.900 17.980 4.140 ;
        RECT  5.390 1.130 18.140 1.370 ;
        RECT  17.680 1.130 18.140 1.550 ;
        RECT  11.820 1.130 12.060 2.900 ;
        RECT  17.900 1.130 18.140 3.550 ;
        RECT  11.960 2.600 12.200 3.570 ;
        RECT  5.390 1.130 5.630 3.650 ;
        RECT  5.170 3.330 5.630 3.650 ;
        RECT  19.270 1.650 19.510 3.580 ;
        RECT  19.270 3.180 21.000 3.580 ;
        RECT  18.450 1.170 19.990 1.410 ;
        RECT  18.450 1.170 18.880 1.900 ;
        RECT  19.750 1.170 19.990 2.460 ;
        RECT  19.750 2.220 21.310 2.460 ;
        RECT  18.640 1.170 18.880 3.550 ;
        RECT  21.160 1.580 21.790 1.980 ;
        RECT  20.230 2.700 21.790 2.940 ;
        RECT  21.550 1.580 21.790 4.140 ;
        RECT  21.550 3.900 22.310 4.140 ;
        RECT  22.220 1.950 22.460 3.470 ;
        RECT  15.270 3.420 15.510 4.370 ;
        RECT  23.210 3.940 23.790 4.180 ;
        RECT  18.700 4.100 21.040 4.340 ;
        RECT  15.270 4.130 17.180 4.370 ;
        RECT  16.940 4.130 17.180 4.620 ;
        RECT  20.800 4.100 21.040 4.620 ;
        RECT  18.700 4.100 18.940 4.620 ;
        RECT  16.940 4.380 18.940 4.620 ;
        RECT  23.210 1.460 23.450 4.620 ;
        RECT  20.800 4.380 23.450 4.620 ;
        RECT  22.030 0.980 23.930 1.220 ;
        RECT  22.030 0.980 22.270 1.710 ;
        RECT  23.690 0.980 23.930 2.720 ;
        RECT  23.690 2.480 24.480 2.720 ;
        RECT  22.730 0.980 22.970 4.140 ;
        RECT  25.030 1.690 25.610 1.930 ;
        RECT  25.370 2.220 25.930 2.460 ;
        RECT  23.720 3.080 23.960 3.700 ;
        RECT  25.370 1.690 25.610 3.700 ;
        RECT  23.720 3.460 25.610 3.700 ;
    END
END secrq2

MACRO secrq1
    CLASS CORE ;
    FOREIGN secrq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.880 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.419  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  24.720 2.400 25.130 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.405  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.720 2.510 16.330 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.940 2.250 13.380 3.020 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.397  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.700 2.580 7.310 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  26.240 3.190 26.740 3.510 ;
        RECT  26.460 1.480 26.740 3.510 ;
        RECT  26.330 1.480 26.740 1.800 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.020 0.980 2.900 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.280 1.640 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 26.880 5.600 ;
        RECT  25.540 4.190 25.780 5.600 ;
        RECT  24.240 4.190 24.480 5.600 ;
        RECT  20.080 4.580 20.480 5.600 ;
        RECT  16.280 4.710 16.680 5.600 ;
        RECT  14.640 4.710 15.040 5.600 ;
        RECT  13.390 4.710 13.790 5.600 ;
        RECT  9.670 4.480 10.070 5.600 ;
        RECT  8.200 3.770 8.440 5.600 ;
        RECT  6.900 3.770 7.140 5.600 ;
        RECT  6.000 3.850 6.240 5.600 ;
        RECT  3.930 4.090 4.170 5.600 ;
        RECT  1.660 4.460 2.060 5.600 ;
        RECT  0.970 3.290 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 26.880 0.740 ;
        RECT  25.670 0.000 25.910 1.300 ;
        RECT  20.470 0.000 20.710 1.980 ;
        RECT  16.460 0.000 16.860 0.890 ;
        RECT  15.050 0.000 15.450 0.890 ;
        RECT  13.070 0.000 13.470 0.890 ;
        RECT  10.170 0.000 10.570 0.890 ;
        RECT  8.130 0.000 8.530 0.890 ;
        RECT  6.180 0.000 6.600 0.890 ;
        RECT  4.190 0.000 4.430 1.470 ;
        RECT  1.660 0.000 2.060 1.140 ;
        RECT  0.760 0.000 1.180 1.180 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 1.520 0.470 1.920 ;
        RECT  0.220 1.520 0.460 4.620 ;
        RECT  0.220 3.290 0.470 4.620 ;
        RECT  1.570 1.530 2.120 1.850 ;
        RECT  1.880 2.270 2.990 2.510 ;
        RECT  1.880 1.530 2.120 3.650 ;
        RECT  1.630 3.330 2.120 3.650 ;
        RECT  2.430 0.980 2.990 1.380 ;
        RECT  2.670 0.980 2.990 1.910 ;
        RECT  2.670 1.630 3.470 1.910 ;
        RECT  3.230 1.630 3.470 2.990 ;
        RECT  2.480 2.750 3.470 2.990 ;
        RECT  2.480 2.750 2.720 4.620 ;
        RECT  2.430 4.220 2.830 4.620 ;
        RECT  3.230 1.150 3.950 1.390 ;
        RECT  3.710 2.800 4.450 3.040 ;
        RECT  3.710 1.150 3.950 3.610 ;
        RECT  2.960 3.370 3.950 3.610 ;
        RECT  2.960 3.370 3.280 3.770 ;
        RECT  4.570 1.830 4.930 2.150 ;
        RECT  4.690 1.830 4.930 3.750 ;
        RECT  4.430 3.430 4.930 3.750 ;
        RECT  6.000 1.610 6.580 1.850 ;
        RECT  6.000 1.610 6.240 3.510 ;
        RECT  9.440 1.610 9.680 2.500 ;
        RECT  9.160 2.260 10.280 2.500 ;
        RECT  9.160 2.260 9.400 3.740 ;
        RECT  10.170 1.690 10.760 1.930 ;
        RECT  10.520 1.690 10.760 3.740 ;
        RECT  10.520 2.510 11.050 2.910 ;
        RECT  10.520 2.510 10.840 3.740 ;
        RECT  10.440 3.340 10.840 3.740 ;
        RECT  12.460 1.610 12.880 1.930 ;
        RECT  12.460 1.610 12.700 3.510 ;
        RECT  12.460 3.270 13.020 3.510 ;
        RECT  6.900 1.620 7.860 1.860 ;
        RECT  7.620 1.620 7.860 3.510 ;
        RECT  7.540 3.110 7.940 3.510 ;
        RECT  7.540 3.270 8.920 3.510 ;
        RECT  8.680 3.270 8.920 4.240 ;
        RECT  8.680 4.000 10.600 4.240 ;
        RECT  10.360 4.000 10.600 4.530 ;
        RECT  12.900 4.230 14.140 4.470 ;
        RECT  10.360 4.290 13.140 4.530 ;
        RECT  13.930 1.610 14.170 2.540 ;
        RECT  13.930 2.140 14.530 2.540 ;
        RECT  14.070 2.140 14.310 3.510 ;
        RECT  11.000 1.610 11.540 1.930 ;
        RECT  14.790 1.630 15.450 2.030 ;
        RECT  11.300 1.610 11.540 4.050 ;
        RECT  11.140 3.250 11.540 4.050 ;
        RECT  12.400 3.750 15.030 3.990 ;
        RECT  11.140 3.810 12.700 4.050 ;
        RECT  14.790 1.630 15.030 4.350 ;
        RECT  15.850 1.910 16.810 2.150 ;
        RECT  16.570 2.760 17.180 3.000 ;
        RECT  16.570 1.910 16.810 3.530 ;
        RECT  15.750 3.290 16.810 3.530 ;
        RECT  17.150 1.830 17.660 2.150 ;
        RECT  17.050 3.290 17.660 3.530 ;
        RECT  17.420 1.830 17.660 4.140 ;
        RECT  17.420 3.900 17.980 4.140 ;
        RECT  5.390 1.130 18.140 1.370 ;
        RECT  17.680 1.130 18.140 1.550 ;
        RECT  11.820 1.130 12.060 2.900 ;
        RECT  17.900 1.130 18.140 3.550 ;
        RECT  11.960 2.600 12.200 3.570 ;
        RECT  5.390 1.130 5.630 3.650 ;
        RECT  5.170 3.330 5.630 3.650 ;
        RECT  19.270 1.650 19.510 3.580 ;
        RECT  19.270 3.180 21.000 3.580 ;
        RECT  18.450 1.170 19.990 1.410 ;
        RECT  18.450 1.170 18.880 1.900 ;
        RECT  19.750 1.170 19.990 2.460 ;
        RECT  19.750 2.220 21.310 2.460 ;
        RECT  18.640 1.170 18.880 3.550 ;
        RECT  21.160 1.660 21.790 1.900 ;
        RECT  20.230 2.700 21.790 2.940 ;
        RECT  21.550 1.660 21.790 4.140 ;
        RECT  21.550 3.900 22.310 4.140 ;
        RECT  22.220 1.950 22.460 3.470 ;
        RECT  15.270 3.420 15.510 4.370 ;
        RECT  23.210 3.940 23.790 4.180 ;
        RECT  18.700 4.100 21.040 4.340 ;
        RECT  15.270 4.130 17.180 4.370 ;
        RECT  16.940 4.130 17.180 4.620 ;
        RECT  20.800 4.100 21.040 4.620 ;
        RECT  18.700 4.100 18.940 4.620 ;
        RECT  16.940 4.380 18.940 4.620 ;
        RECT  23.210 1.460 23.450 4.620 ;
        RECT  20.800 4.380 23.450 4.620 ;
        RECT  22.030 0.980 23.930 1.220 ;
        RECT  22.030 0.980 22.270 1.710 ;
        RECT  23.690 0.980 23.930 2.720 ;
        RECT  23.690 2.480 24.480 2.720 ;
        RECT  22.730 0.980 22.970 4.140 ;
        RECT  25.060 1.690 25.610 1.930 ;
        RECT  25.370 2.220 25.930 2.460 ;
        RECT  23.720 3.080 23.960 3.700 ;
        RECT  25.370 1.690 25.610 3.700 ;
        RECT  23.720 3.460 25.610 3.700 ;
    END
END secrq1

MACRO secfq4
    CLASS CORE ;
    FOREIGN secfq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.440 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.949  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.710 2.420 12.260 3.020 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.515  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  26.940 2.300 27.320 3.020 ;
        RECT  26.640 2.300 27.320 2.700 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.710 2.040 2.180 2.440 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.510 0.570 3.020 ;
        RECT  0.170 2.410 0.570 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.092  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  23.700 2.940 24.280 3.180 ;
        RECT  20.940 3.010 23.810 3.200 ;
        RECT  21.370 2.960 24.280 3.180 ;
        RECT  23.020 2.580 23.460 3.200 ;
        RECT  23.040 1.560 23.360 3.200 ;
        RECT  21.560 1.880 23.360 2.120 ;
        RECT  22.960 1.560 23.360 2.120 ;
        RECT  21.560 1.460 21.800 2.120 ;
        RECT  20.940 3.010 21.580 3.250 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.531  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.130 2.580 7.780 3.020 ;
        RECT  7.130 2.330 7.530 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.362  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.280 3.140 6.100 3.580 ;
        RECT  5.280 2.120 5.700 3.580 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 27.440 5.600 ;
        RECT  26.380 4.450 26.620 5.600 ;
        RECT  25.680 3.170 25.920 5.600 ;
        RECT  24.290 4.410 24.530 5.600 ;
        RECT  23.180 4.350 23.420 5.600 ;
        RECT  21.730 4.050 21.970 5.600 ;
        RECT  20.280 4.310 20.520 5.600 ;
        RECT  19.000 4.020 19.240 5.600 ;
        RECT  14.360 4.400 14.600 5.600 ;
        RECT  12.880 4.400 13.120 5.600 ;
        RECT  11.440 4.400 11.680 5.600 ;
        RECT  7.920 4.450 8.160 5.600 ;
        RECT  6.470 4.300 6.710 5.600 ;
        RECT  3.320 4.050 3.560 5.600 ;
        RECT  0.230 4.250 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 27.440 0.740 ;
        RECT  25.880 0.000 26.120 1.570 ;
        RECT  23.810 0.000 24.050 1.260 ;
        RECT  22.300 0.000 22.540 1.640 ;
        RECT  20.820 0.000 21.060 1.640 ;
        RECT  16.510 0.000 16.750 1.700 ;
        RECT  13.540 0.000 13.780 1.260 ;
        RECT  8.130 0.000 8.530 0.900 ;
        RECT  5.460 0.000 5.860 0.900 ;
        RECT  2.770 0.000 3.170 0.890 ;
        RECT  0.150 0.000 0.550 0.960 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 2.420 1.330 2.820 ;
        RECT  4.150 2.590 4.550 2.990 ;
        RECT  0.820 1.670 1.060 3.990 ;
        RECT  2.280 3.510 4.390 3.750 ;
        RECT  4.150 2.590 4.390 3.750 ;
        RECT  0.820 3.750 2.520 3.990 ;
        RECT  3.030 1.140 6.360 1.380 ;
        RECT  6.120 1.620 7.460 1.860 ;
        RECT  3.030 1.140 3.270 2.450 ;
        RECT  7.220 1.850 8.010 2.090 ;
        RECT  7.770 2.260 8.330 2.340 ;
        RECT  7.770 1.850 8.010 2.340 ;
        RECT  3.030 2.030 3.430 2.450 ;
        RECT  8.010 2.290 8.360 2.500 ;
        RECT  8.010 2.090 8.240 2.500 ;
        RECT  5.990 2.500 6.390 2.900 ;
        RECT  8.120 2.490 8.520 2.890 ;
        RECT  6.120 1.140 6.360 2.900 ;
        RECT  6.340 2.660 6.580 3.580 ;
        RECT  6.340 3.340 7.590 3.580 ;
        RECT  6.600 0.980 7.000 1.380 ;
        RECT  6.600 1.140 8.030 1.380 ;
        RECT  7.790 1.360 8.810 1.600 ;
        RECT  8.510 1.360 8.810 2.100 ;
        RECT  8.510 1.700 9.180 2.100 ;
        RECT  8.940 1.700 9.180 3.370 ;
        RECT  8.520 3.130 9.180 3.370 ;
        RECT  9.110 0.980 9.660 1.220 ;
        RECT  1.540 1.540 2.660 1.780 ;
        RECT  4.790 1.620 5.420 1.860 ;
        RECT  3.670 1.860 5.030 2.100 ;
        RECT  2.420 2.690 3.910 2.930 ;
        RECT  3.670 1.860 3.910 2.930 ;
        RECT  2.420 1.540 2.660 2.940 ;
        RECT  1.760 2.700 2.660 2.940 ;
        RECT  1.760 2.700 2.000 3.510 ;
        RECT  1.440 3.270 2.000 3.510 ;
        RECT  4.790 1.620 5.030 4.060 ;
        RECT  4.790 3.820 8.990 4.060 ;
        RECT  9.420 0.980 9.660 4.620 ;
        RECT  8.750 3.820 8.990 4.540 ;
        RECT  5.050 3.820 5.450 4.310 ;
        RECT  8.750 4.300 9.680 4.540 ;
        RECT  9.280 4.220 9.680 4.620 ;
        RECT  10.720 1.510 10.960 2.390 ;
        RECT  10.410 2.150 10.960 2.390 ;
        RECT  10.410 2.150 10.650 3.270 ;
        RECT  10.410 3.030 10.900 3.270 ;
        RECT  10.660 3.030 10.900 4.620 ;
        RECT  10.660 3.920 12.160 4.160 ;
        RECT  11.920 3.920 12.160 4.620 ;
        RECT  10.610 4.160 11.010 4.620 ;
        RECT  11.920 4.380 12.500 4.620 ;
        RECT  9.900 0.980 12.040 1.220 ;
        RECT  11.800 0.980 12.040 1.520 ;
        RECT  11.800 1.280 13.290 1.520 ;
        RECT  13.050 1.510 14.010 1.750 ;
        RECT  9.900 1.510 10.300 1.910 ;
        RECT  13.560 1.510 14.010 1.910 ;
        RECT  9.900 0.980 10.140 3.920 ;
        RECT  9.900 3.520 10.420 3.920 ;
        RECT  14.300 1.320 16.130 1.560 ;
        RECT  15.730 1.290 16.130 1.700 ;
        RECT  12.560 1.760 12.800 2.390 ;
        RECT  14.300 1.320 14.540 2.390 ;
        RECT  12.560 2.150 14.540 2.390 ;
        RECT  17.470 1.980 17.710 2.660 ;
        RECT  15.410 2.420 17.710 2.660 ;
        RECT  15.410 2.420 15.650 3.370 ;
        RECT  15.170 3.130 15.650 3.370 ;
        RECT  11.140 2.820 11.380 3.680 ;
        RECT  11.140 3.440 12.650 3.680 ;
        RECT  12.410 3.440 12.650 4.000 ;
        RECT  12.410 3.760 15.420 4.000 ;
        RECT  15.180 3.950 16.300 4.190 ;
        RECT  15.180 3.130 15.420 4.620 ;
        RECT  18.240 1.550 18.480 2.130 ;
        RECT  18.190 1.890 18.430 3.140 ;
        RECT  15.910 2.900 18.430 3.140 ;
        RECT  15.910 2.900 16.310 3.300 ;
        RECT  17.430 2.900 17.670 4.010 ;
        RECT  17.430 3.610 17.960 4.010 ;
        RECT  16.990 0.980 20.580 1.220 ;
        RECT  14.810 1.880 15.570 2.120 ;
        RECT  16.990 0.980 17.230 2.180 ;
        RECT  15.400 1.940 17.230 2.180 ;
        RECT  20.340 0.980 20.580 2.710 ;
        RECT  19.980 2.300 21.130 2.710 ;
        RECT  19.980 2.360 22.750 2.710 ;
        RECT  14.810 1.880 15.050 2.870 ;
        RECT  13.620 2.630 15.050 2.870 ;
        RECT  19.980 2.300 20.220 3.290 ;
        RECT  19.820 2.890 20.220 3.290 ;
        RECT  13.620 2.630 13.860 3.520 ;
        RECT  24.700 0.980 25.100 1.380 ;
        RECT  24.400 1.140 25.100 1.380 ;
        RECT  18.900 1.460 19.300 1.860 ;
        RECT  18.900 1.620 20.100 1.860 ;
        RECT  18.900 1.460 19.140 2.610 ;
        RECT  24.400 1.140 24.640 2.610 ;
        RECT  18.670 2.370 18.910 3.780 ;
        RECT  23.100 3.440 24.770 3.680 ;
        RECT  24.530 2.370 24.770 3.680 ;
        RECT  18.460 3.540 20.060 3.780 ;
        RECT  19.660 3.570 23.340 3.810 ;
        RECT  19.660 3.540 20.060 4.020 ;
        RECT  18.460 3.540 18.700 4.610 ;
        RECT  18.150 4.370 18.700 4.610 ;
        RECT  24.900 1.620 25.310 2.020 ;
        RECT  25.070 1.620 25.310 4.170 ;
        RECT  23.660 3.930 25.330 4.170 ;
        RECT  23.660 3.930 24.060 4.330 ;
        RECT  25.090 3.930 25.330 4.580 ;
        RECT  26.540 1.580 26.940 2.050 ;
        RECT  25.770 1.810 26.940 2.050 ;
        RECT  25.770 1.810 26.010 2.920 ;
        RECT  25.750 2.520 26.170 2.920 ;
        RECT  26.160 2.550 26.400 3.510 ;
        RECT  26.160 3.270 27.290 3.510 ;
    END
END secfq4

MACRO secfq2
    CLASS CORE ;
    FOREIGN secfq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.760 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.941  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.710 2.420 12.260 3.020 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.515  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  25.260 2.480 25.640 3.020 ;
        RECT  24.720 2.480 25.640 2.880 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.710 2.040 2.180 2.440 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.510 0.570 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.394  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  20.940 3.340 21.800 3.580 ;
        RECT  21.560 1.460 21.800 3.580 ;
        RECT  21.340 2.580 21.800 3.580 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.419  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.110 2.580 7.780 3.020 ;
        RECT  7.110 2.330 7.510 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.280 3.140 6.100 3.580 ;
        RECT  5.280 2.120 5.700 3.580 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 25.760 5.600 ;
        RECT  24.700 4.450 24.940 5.600 ;
        RECT  23.500 4.260 23.740 5.600 ;
        RECT  23.180 4.260 23.740 4.500 ;
        RECT  21.580 4.350 21.820 5.600 ;
        RECT  20.280 4.310 20.520 5.600 ;
        RECT  19.000 4.020 19.240 5.600 ;
        RECT  14.440 4.400 14.680 5.600 ;
        RECT  12.880 4.400 13.120 5.600 ;
        RECT  11.440 4.400 11.680 5.600 ;
        RECT  7.640 4.300 8.240 4.540 ;
        RECT  7.640 4.300 7.880 5.600 ;
        RECT  6.470 4.310 6.710 5.600 ;
        RECT  3.320 4.050 3.560 5.600 ;
        RECT  0.230 4.250 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 25.760 0.740 ;
        RECT  24.390 0.000 24.630 1.510 ;
        RECT  22.330 0.000 22.570 1.270 ;
        RECT  20.820 0.000 21.060 1.640 ;
        RECT  16.510 0.000 16.750 1.700 ;
        RECT  13.540 0.000 13.780 1.260 ;
        RECT  8.130 0.000 8.530 0.900 ;
        RECT  5.460 0.000 5.860 0.900 ;
        RECT  2.770 0.000 3.170 0.890 ;
        RECT  0.150 0.000 0.550 1.060 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 2.520 1.330 2.920 ;
        RECT  4.150 2.590 4.550 2.990 ;
        RECT  0.820 1.770 1.060 3.990 ;
        RECT  2.280 3.510 4.390 3.750 ;
        RECT  4.150 2.590 4.390 3.750 ;
        RECT  0.820 3.750 2.520 3.990 ;
        RECT  3.030 1.140 6.360 1.380 ;
        RECT  6.120 1.650 7.460 1.890 ;
        RECT  3.030 1.140 3.270 2.450 ;
        RECT  7.220 1.850 8.010 2.090 ;
        RECT  7.770 2.260 8.330 2.340 ;
        RECT  7.770 1.850 8.010 2.340 ;
        RECT  3.030 2.030 3.430 2.450 ;
        RECT  8.010 2.290 8.360 2.500 ;
        RECT  8.010 2.090 8.240 2.500 ;
        RECT  5.990 2.500 6.390 2.900 ;
        RECT  8.120 2.490 8.520 2.890 ;
        RECT  6.120 1.140 6.360 2.900 ;
        RECT  6.340 2.660 6.580 3.580 ;
        RECT  6.340 3.340 7.590 3.580 ;
        RECT  6.600 1.010 7.000 1.410 ;
        RECT  6.600 1.120 8.030 1.410 ;
        RECT  7.790 1.360 8.810 1.600 ;
        RECT  8.510 1.360 8.810 2.100 ;
        RECT  8.510 1.700 9.180 2.100 ;
        RECT  8.940 1.700 9.180 3.370 ;
        RECT  8.520 3.130 9.180 3.370 ;
        RECT  9.110 0.980 9.660 1.220 ;
        RECT  1.540 1.540 2.660 1.780 ;
        RECT  4.790 1.620 5.420 1.860 ;
        RECT  3.670 1.860 5.030 2.100 ;
        RECT  2.420 2.690 3.910 2.930 ;
        RECT  3.670 1.860 3.910 2.930 ;
        RECT  2.420 1.540 2.660 2.940 ;
        RECT  1.760 2.700 2.660 2.940 ;
        RECT  1.760 2.700 2.000 3.510 ;
        RECT  1.440 3.270 2.000 3.510 ;
        RECT  4.790 1.620 5.030 4.060 ;
        RECT  4.790 3.820 8.990 4.060 ;
        RECT  9.420 0.980 9.660 4.620 ;
        RECT  8.750 3.820 8.990 4.540 ;
        RECT  5.050 3.820 5.450 4.310 ;
        RECT  8.750 4.300 9.680 4.540 ;
        RECT  9.280 4.220 9.680 4.620 ;
        RECT  10.700 1.510 10.940 2.390 ;
        RECT  10.660 2.150 10.900 4.620 ;
        RECT  10.660 3.920 12.160 4.160 ;
        RECT  11.920 3.920 12.160 4.620 ;
        RECT  10.610 4.160 11.010 4.620 ;
        RECT  11.920 4.380 12.500 4.620 ;
        RECT  9.960 0.980 12.040 1.220 ;
        RECT  11.800 0.980 12.040 1.520 ;
        RECT  11.800 1.280 13.290 1.520 ;
        RECT  13.050 1.510 14.010 1.750 ;
        RECT  13.560 1.510 14.010 1.910 ;
        RECT  9.960 0.980 10.200 3.920 ;
        RECT  9.960 3.520 10.420 3.920 ;
        RECT  14.300 1.290 16.130 1.530 ;
        RECT  15.730 1.290 16.130 1.700 ;
        RECT  12.560 1.760 12.800 2.390 ;
        RECT  14.300 1.290 14.540 2.390 ;
        RECT  12.560 2.150 14.540 2.390 ;
        RECT  17.470 1.980 17.790 2.660 ;
        RECT  15.410 2.420 17.790 2.660 ;
        RECT  15.410 2.420 15.650 3.370 ;
        RECT  15.170 3.130 15.650 3.370 ;
        RECT  11.140 2.820 11.380 3.680 ;
        RECT  11.140 3.440 12.650 3.680 ;
        RECT  12.410 3.440 12.650 4.140 ;
        RECT  12.410 3.900 15.420 4.140 ;
        RECT  15.180 3.950 16.300 4.190 ;
        RECT  15.180 3.130 15.420 4.620 ;
        RECT  18.240 1.550 18.480 2.130 ;
        RECT  18.190 1.890 18.430 3.140 ;
        RECT  15.910 2.900 18.430 3.140 ;
        RECT  15.910 2.900 16.310 3.300 ;
        RECT  17.430 2.900 17.670 4.010 ;
        RECT  17.430 3.610 17.960 4.010 ;
        RECT  16.990 0.980 20.580 1.220 ;
        RECT  14.880 1.770 15.360 2.180 ;
        RECT  16.990 0.980 17.230 2.180 ;
        RECT  14.880 1.940 17.230 2.180 ;
        RECT  20.340 0.980 20.580 2.530 ;
        RECT  19.980 2.290 20.580 2.530 ;
        RECT  14.880 1.770 15.170 2.870 ;
        RECT  13.620 2.630 15.170 2.870 ;
        RECT  19.980 2.290 20.220 3.300 ;
        RECT  19.820 2.900 20.220 3.300 ;
        RECT  13.620 2.630 13.860 3.500 ;
        RECT  22.810 1.060 23.610 1.300 ;
        RECT  22.810 1.060 23.050 1.750 ;
        RECT  22.040 1.510 23.050 1.750 ;
        RECT  18.900 1.540 20.100 1.790 ;
        RECT  19.700 1.540 20.100 1.940 ;
        RECT  18.900 1.540 19.300 2.610 ;
        RECT  18.670 2.370 18.910 3.780 ;
        RECT  18.460 3.540 20.060 3.780 ;
        RECT  19.660 3.540 20.060 4.070 ;
        RECT  22.040 1.510 22.280 4.070 ;
        RECT  19.660 3.830 22.280 4.070 ;
        RECT  18.460 3.540 18.700 4.610 ;
        RECT  18.150 4.370 18.700 4.610 ;
        RECT  23.290 1.590 23.850 1.830 ;
        RECT  23.290 1.590 23.530 2.730 ;
        RECT  22.620 2.490 23.530 2.730 ;
        RECT  22.620 2.490 23.030 2.890 ;
        RECT  22.790 2.490 23.030 3.960 ;
        RECT  22.520 3.720 24.320 3.960 ;
        RECT  22.520 3.720 22.760 4.290 ;
        RECT  25.050 1.520 25.450 2.010 ;
        RECT  24.110 1.770 25.450 2.010 ;
        RECT  24.110 1.770 24.350 3.370 ;
        RECT  23.430 3.130 24.800 3.370 ;
        RECT  23.430 3.060 23.830 3.460 ;
        RECT  24.560 3.270 25.610 3.510 ;
    END
END secfq2

MACRO secfq1
    CLASS CORE ;
    FOREIGN secfq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.950  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.710 2.420 12.260 3.020 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.504  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  23.580 2.580 24.020 3.020 ;
        RECT  23.330 2.560 23.730 2.960 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.710 2.040 2.180 2.440 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.510 0.570 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.160  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  21.450 1.070 22.060 1.310 ;
        RECT  20.970 1.900 21.690 2.140 ;
        RECT  21.450 1.070 21.690 2.140 ;
        RECT  20.340 2.840 21.210 3.080 ;
        RECT  20.970 1.900 21.210 3.080 ;
        RECT  20.220 3.180 20.740 3.580 ;
        RECT  20.340 2.840 20.740 3.580 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.531  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.210 2.580 7.780 3.020 ;
        RECT  7.210 2.330 7.610 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.362  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.280 3.140 6.100 3.580 ;
        RECT  5.280 2.120 5.700 3.580 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 24.640 5.600 ;
        RECT  22.820 4.440 23.060 5.600 ;
        RECT  18.970 3.860 19.210 5.600 ;
        RECT  14.440 4.400 14.680 5.600 ;
        RECT  12.880 4.400 13.120 5.600 ;
        RECT  11.440 4.400 11.680 5.600 ;
        RECT  7.780 4.610 8.180 5.600 ;
        RECT  6.470 4.300 6.710 5.600 ;
        RECT  3.320 4.050 3.560 5.600 ;
        RECT  0.230 4.250 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 24.640 0.740 ;
        RECT  23.000 0.000 23.400 0.890 ;
        RECT  20.970 0.000 21.210 1.660 ;
        RECT  16.660 0.000 16.900 1.700 ;
        RECT  13.650 0.000 13.890 1.260 ;
        RECT  8.130 0.000 8.530 0.900 ;
        RECT  5.460 0.000 5.860 0.900 ;
        RECT  2.770 0.000 3.170 0.890 ;
        RECT  0.150 0.000 0.550 1.060 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 2.520 1.330 2.920 ;
        RECT  4.150 2.590 4.550 2.990 ;
        RECT  0.820 1.770 1.060 3.990 ;
        RECT  2.280 3.510 4.390 3.750 ;
        RECT  4.150 2.590 4.390 3.750 ;
        RECT  0.820 3.750 2.520 3.990 ;
        RECT  3.030 1.140 6.360 1.380 ;
        RECT  6.120 1.620 7.460 1.860 ;
        RECT  3.030 1.140 3.270 2.450 ;
        RECT  7.220 1.850 8.250 2.090 ;
        RECT  3.030 2.030 3.430 2.450 ;
        RECT  8.010 1.850 8.250 2.510 ;
        RECT  5.990 2.500 6.390 2.900 ;
        RECT  8.020 2.440 8.520 2.890 ;
        RECT  6.120 1.140 6.360 2.900 ;
        RECT  6.340 2.660 6.580 3.580 ;
        RECT  6.340 3.340 7.590 3.580 ;
        RECT  6.600 0.980 7.000 1.380 ;
        RECT  6.600 1.140 8.030 1.380 ;
        RECT  7.790 1.360 8.730 1.600 ;
        RECT  8.490 1.360 8.730 2.100 ;
        RECT  8.490 1.700 8.890 2.100 ;
        RECT  8.490 1.860 9.180 2.100 ;
        RECT  8.940 1.860 9.180 3.370 ;
        RECT  8.520 3.130 9.180 3.370 ;
        RECT  9.110 0.980 9.660 1.220 ;
        RECT  1.540 1.540 2.660 1.780 ;
        RECT  4.790 1.620 5.420 1.860 ;
        RECT  3.670 1.860 5.030 2.100 ;
        RECT  2.420 2.690 3.910 2.930 ;
        RECT  3.670 1.860 3.910 2.930 ;
        RECT  2.420 1.540 2.660 2.940 ;
        RECT  1.760 2.700 2.660 2.940 ;
        RECT  1.760 2.700 2.000 3.510 ;
        RECT  1.440 3.270 2.000 3.510 ;
        RECT  4.790 1.620 5.030 4.060 ;
        RECT  4.790 3.820 7.190 4.060 ;
        RECT  6.950 3.820 7.190 4.360 ;
        RECT  9.420 0.980 9.660 4.620 ;
        RECT  5.050 3.820 5.450 4.310 ;
        RECT  6.950 4.120 8.660 4.360 ;
        RECT  8.420 4.300 9.680 4.540 ;
        RECT  9.280 4.220 9.680 4.620 ;
        RECT  10.700 1.510 10.940 2.390 ;
        RECT  10.660 2.150 10.900 4.620 ;
        RECT  10.660 3.920 12.160 4.160 ;
        RECT  11.920 3.920 12.160 4.620 ;
        RECT  10.610 4.160 11.010 4.620 ;
        RECT  11.920 4.380 12.500 4.620 ;
        RECT  9.960 0.980 12.040 1.220 ;
        RECT  11.800 0.980 12.040 1.520 ;
        RECT  11.800 1.280 13.410 1.520 ;
        RECT  13.170 1.510 14.110 1.750 ;
        RECT  13.710 1.510 14.110 1.910 ;
        RECT  9.960 0.980 10.200 3.920 ;
        RECT  9.960 3.520 10.420 3.920 ;
        RECT  14.450 1.290 16.280 1.530 ;
        RECT  15.880 1.290 16.280 1.700 ;
        RECT  12.670 1.760 12.910 2.390 ;
        RECT  14.450 1.290 14.690 2.390 ;
        RECT  12.670 2.150 14.690 2.390 ;
        RECT  17.620 1.980 17.860 2.660 ;
        RECT  15.410 2.420 17.860 2.660 ;
        RECT  15.410 2.420 15.650 3.370 ;
        RECT  15.170 3.130 15.650 3.370 ;
        RECT  11.140 2.820 11.380 3.680 ;
        RECT  11.140 3.440 12.650 3.680 ;
        RECT  12.410 3.440 12.650 4.140 ;
        RECT  12.410 3.900 15.420 4.140 ;
        RECT  15.180 3.950 16.300 4.190 ;
        RECT  15.180 3.130 15.420 4.620 ;
        RECT  18.390 1.550 18.630 2.130 ;
        RECT  18.190 1.890 18.430 3.140 ;
        RECT  15.910 2.900 18.430 3.140 ;
        RECT  15.910 2.900 16.310 3.300 ;
        RECT  17.430 2.900 17.670 4.010 ;
        RECT  17.430 3.610 17.960 4.010 ;
        RECT  17.140 0.980 20.730 1.220 ;
        RECT  14.930 1.770 15.510 2.180 ;
        RECT  17.140 0.980 17.380 2.180 ;
        RECT  14.930 1.940 17.380 2.180 ;
        RECT  20.490 0.980 20.730 2.530 ;
        RECT  19.850 2.290 20.730 2.530 ;
        RECT  14.930 1.770 15.170 2.870 ;
        RECT  13.670 2.630 15.170 2.870 ;
        RECT  19.850 2.290 20.090 2.950 ;
        RECT  19.680 2.550 20.090 2.950 ;
        RECT  13.670 2.630 13.910 3.500 ;
        RECT  21.930 1.730 22.630 1.970 ;
        RECT  21.930 1.730 22.170 2.710 ;
        RECT  21.480 2.470 22.090 2.870 ;
        RECT  21.850 2.470 22.090 3.770 ;
        RECT  22.870 1.640 23.990 1.880 ;
        RECT  22.870 1.640 23.110 2.450 ;
        RECT  22.410 2.210 23.110 2.450 ;
        RECT  22.410 2.210 22.810 2.610 ;
        RECT  22.570 2.210 22.810 3.500 ;
        RECT  22.570 3.260 23.890 3.500 ;
        RECT  23.950 0.980 24.500 1.380 ;
        RECT  19.050 1.550 20.250 1.790 ;
        RECT  19.050 1.550 19.450 1.950 ;
        RECT  19.850 1.550 20.250 2.050 ;
        RECT  19.050 1.550 19.340 2.610 ;
        RECT  18.670 2.370 19.340 2.610 ;
        RECT  18.670 2.370 18.910 3.620 ;
        RECT  18.460 3.380 19.710 3.620 ;
        RECT  19.470 3.380 19.710 4.190 ;
        RECT  19.470 3.950 21.680 4.190 ;
        RECT  22.260 3.950 24.500 4.190 ;
        RECT  24.260 0.980 24.500 4.190 ;
        RECT  18.460 3.380 18.700 4.610 ;
        RECT  21.440 4.190 22.500 4.430 ;
        RECT  18.150 4.370 18.700 4.610 ;
    END
END secfq1

MACRO sdprb4
    CLASS CORE ;
    FOREIGN sdprb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.000 5.620 2.460 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.020 2.740 2.460 ;
        RECT  2.480 1.620 2.720 2.460 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.881  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  20.780 1.460 21.160 1.900 ;
        RECT  18.400 1.460 21.160 1.700 ;
        RECT  18.630 3.350 20.340 3.590 ;
        RECT  19.070 1.460 19.310 3.590 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.036  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.980 2.580 18.420 3.020 ;
        RECT  16.220 1.460 18.100 1.700 ;
        RECT  17.400 2.580 18.420 2.820 ;
        RECT  17.320 3.600 17.720 4.000 ;
        RECT  17.400 1.460 17.640 4.000 ;
        RECT  15.960 3.680 17.720 3.920 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.480 2.030 0.720 2.820 ;
        RECT  0.120 2.580 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.020 4.410 3.080 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.794  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.700 2.420 14.940 3.990 ;
        RECT  13.390 3.750 14.940 3.990 ;
        RECT  13.140 2.420 14.940 2.660 ;
        RECT  10.940 3.960 13.630 4.200 ;
        RECT  12.940 2.020 13.380 2.460 ;
        RECT  10.940 2.390 11.180 4.200 ;
        RECT  9.690 2.390 11.180 2.630 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 21.280 5.600 ;
        RECT  20.680 4.620 21.080 5.600 ;
        RECT  19.370 4.620 19.770 5.600 ;
        RECT  18.060 4.620 18.460 5.600 ;
        RECT  16.760 4.620 17.160 5.600 ;
        RECT  15.430 4.710 15.830 5.600 ;
        RECT  13.270 4.710 13.670 5.600 ;
        RECT  10.290 4.710 10.690 5.600 ;
        RECT  8.880 4.710 9.280 5.600 ;
        RECT  5.520 4.330 5.920 5.600 ;
        RECT  3.200 4.380 3.600 5.600 ;
        RECT  0.720 4.400 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 21.280 0.740 ;
        RECT  20.650 0.000 21.050 1.220 ;
        RECT  19.170 0.000 19.570 1.220 ;
        RECT  16.960 0.000 17.360 1.220 ;
        RECT  15.450 0.000 15.850 0.890 ;
        RECT  13.550 0.000 13.950 0.890 ;
        RECT  9.470 1.360 10.370 1.600 ;
        RECT  10.130 0.000 10.370 1.600 ;
        RECT  5.780 0.000 6.180 0.890 ;
        RECT  3.440 0.000 3.840 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.310 1.200 1.550 ;
        RECT  0.960 2.110 1.500 2.510 ;
        RECT  0.960 1.310 1.200 3.510 ;
        RECT  0.150 3.270 1.200 3.510 ;
        RECT  1.510 1.470 1.980 1.870 ;
        RECT  1.740 1.470 1.980 3.110 ;
        RECT  3.020 2.310 3.260 3.110 ;
        RECT  1.510 2.870 3.260 3.110 ;
        RECT  1.510 2.870 1.750 4.610 ;
        RECT  1.460 4.210 1.860 4.610 ;
        RECT  5.190 1.310 6.270 1.550 ;
        RECT  6.030 1.310 6.270 2.940 ;
        RECT  5.950 2.460 6.350 2.940 ;
        RECT  5.050 2.700 6.350 2.940 ;
        RECT  5.050 2.700 5.290 3.480 ;
        RECT  6.550 1.470 7.080 1.870 ;
        RECT  6.840 1.470 7.080 3.420 ;
        RECT  6.270 3.180 7.080 3.420 ;
        RECT  2.210 0.980 3.200 1.220 ;
        RECT  2.960 0.980 3.200 1.760 ;
        RECT  2.960 1.520 4.890 1.760 ;
        RECT  3.500 1.520 3.740 3.600 ;
        RECT  1.990 3.360 4.810 3.600 ;
        RECT  4.570 3.360 4.810 4.080 ;
        RECT  7.330 1.310 7.570 4.080 ;
        RECT  4.570 3.840 7.570 4.080 ;
        RECT  6.880 3.840 7.120 4.620 ;
        RECT  8.630 1.280 9.130 1.680 ;
        RECT  8.630 1.280 8.870 2.110 ;
        RECT  8.300 1.870 8.870 2.110 ;
        RECT  8.300 1.870 8.540 3.450 ;
        RECT  8.300 3.050 8.720 3.450 ;
        RECT  7.810 1.390 8.390 1.630 ;
        RECT  7.810 1.390 8.050 3.980 ;
        RECT  7.810 3.740 8.480 3.980 ;
        RECT  8.240 4.230 10.700 4.470 ;
        RECT  10.460 2.950 10.700 4.470 ;
        RECT  8.240 3.740 8.480 4.610 ;
        RECT  7.540 4.370 8.480 4.610 ;
        RECT  10.750 1.280 10.990 2.150 ;
        RECT  9.210 1.910 11.660 2.150 ;
        RECT  9.210 1.910 9.450 2.590 ;
        RECT  8.780 2.350 9.450 2.590 ;
        RECT  8.780 2.350 9.200 2.750 ;
        RECT  8.960 2.350 9.200 3.880 ;
        RECT  11.420 1.910 11.660 3.720 ;
        RECT  8.960 3.640 10.060 3.880 ;
        RECT  12.380 1.460 12.620 3.140 ;
        RECT  12.380 2.900 14.450 3.140 ;
        RECT  14.210 2.900 14.450 3.510 ;
        RECT  12.910 2.900 13.150 3.720 ;
        RECT  11.900 0.980 13.310 1.220 ;
        RECT  13.070 0.980 13.310 1.780 ;
        RECT  11.410 1.360 12.140 1.600 ;
        RECT  13.070 1.540 13.860 1.780 ;
        RECT  13.620 1.540 13.860 2.180 ;
        RECT  13.620 1.940 15.420 2.180 ;
        RECT  15.180 1.940 15.420 2.800 ;
        RECT  15.180 2.560 16.560 2.800 ;
        RECT  11.900 0.980 12.140 3.640 ;
        RECT  11.900 3.400 12.480 3.640 ;
        RECT  14.120 1.310 15.900 1.550 ;
        RECT  15.660 1.310 15.900 2.180 ;
        RECT  15.660 1.940 17.040 2.180 ;
        RECT  16.800 1.940 17.040 3.440 ;
        RECT  15.180 3.200 17.040 3.440 ;
        RECT  15.180 3.200 15.420 4.470 ;
        RECT  14.660 4.230 15.420 4.470 ;
    END
END sdprb4

MACRO sdprb2
    CLASS CORE ;
    FOREIGN sdprb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.296  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.580 7.630 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.257  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.460 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.420 3.390 20.020 3.630 ;
        RECT  19.740 1.370 20.020 3.630 ;
        RECT  19.420 1.370 20.020 1.610 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.500 3.390 18.340 3.630 ;
        RECT  17.500 1.370 18.340 1.610 ;
        RECT  17.500 1.370 17.780 3.630 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.520 0.460 2.460 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.090  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.550 4.120 6.020 4.520 ;
        RECT  5.740 3.700 6.020 4.520 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.460 2.480 13.100 2.720 ;
        RECT  12.460 2.020 12.820 2.720 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.720 5.600 ;
        RECT  20.240 4.390 20.480 5.600 ;
        RECT  18.760 4.390 19.000 5.600 ;
        RECT  17.280 4.390 17.520 5.600 ;
        RECT  15.280 4.020 15.520 5.600 ;
        RECT  12.480 4.380 12.720 5.600 ;
        RECT  11.130 4.380 11.370 5.600 ;
        RECT  7.220 4.560 7.620 5.600 ;
        RECT  6.180 4.710 6.580 5.600 ;
        RECT  4.870 3.130 5.110 5.600 ;
        RECT  1.900 4.660 2.300 5.600 ;
        RECT  0.430 4.570 0.830 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.720 0.740 ;
        RECT  20.160 0.000 20.560 1.030 ;
        RECT  18.680 0.000 19.080 1.030 ;
        RECT  17.200 0.000 17.600 1.030 ;
        RECT  15.760 0.000 16.160 1.640 ;
        RECT  11.470 0.000 11.710 1.970 ;
        RECT  7.570 0.000 7.970 0.900 ;
        RECT  6.180 0.000 6.580 0.900 ;
        RECT  4.610 0.000 5.010 0.900 ;
        RECT  1.900 0.000 2.300 0.990 ;
        RECT  1.180 0.000 1.420 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.040 0.940 1.280 ;
        RECT  0.700 1.040 0.940 4.230 ;
        RECT  0.430 3.910 0.940 4.230 ;
        RECT  2.540 1.750 2.940 2.070 ;
        RECT  2.700 1.750 2.940 3.690 ;
        RECT  2.540 3.370 2.940 3.690 ;
        RECT  1.210 1.750 1.450 4.230 ;
        RECT  1.210 3.990 3.430 4.230 ;
        RECT  3.030 3.990 3.430 4.390 ;
        RECT  4.020 1.750 4.420 2.070 ;
        RECT  4.020 1.750 4.260 3.690 ;
        RECT  4.020 3.370 4.420 3.690 ;
        RECT  5.350 1.690 5.880 2.010 ;
        RECT  4.510 2.380 5.590 2.620 ;
        RECT  5.350 1.690 5.590 3.370 ;
        RECT  5.350 3.130 5.930 3.370 ;
        RECT  5.870 2.370 6.500 2.610 ;
        RECT  6.260 1.620 6.500 4.370 ;
        RECT  3.360 1.140 9.360 1.380 ;
        RECT  8.870 1.140 9.360 1.640 ;
        RECT  9.060 1.140 9.360 3.600 ;
        RECT  3.360 1.140 3.600 3.690 ;
        RECT  8.360 1.920 8.660 4.140 ;
        RECT  8.360 3.900 9.630 4.140 ;
        RECT  10.350 1.580 10.750 1.980 ;
        RECT  10.460 1.580 10.700 3.600 ;
        RECT  10.460 3.280 10.860 3.600 ;
        RECT  9.610 1.100 11.230 1.340 ;
        RECT  9.610 1.100 10.040 1.850 ;
        RECT  10.990 1.100 11.230 2.450 ;
        RECT  10.990 2.210 12.220 2.450 ;
        RECT  11.980 2.210 12.220 2.800 ;
        RECT  9.800 1.100 10.040 3.600 ;
        RECT  13.030 1.580 13.580 1.900 ;
        RECT  10.950 2.720 11.540 2.960 ;
        RECT  11.300 2.720 11.540 3.600 ;
        RECT  13.340 1.580 13.580 3.600 ;
        RECT  11.300 3.200 13.580 3.600 ;
        RECT  6.980 1.920 8.110 2.160 ;
        RECT  6.980 3.280 8.110 3.520 ;
        RECT  10.400 3.900 13.880 4.140 ;
        RECT  7.870 1.920 8.110 4.620 ;
        RECT  13.640 3.900 13.880 4.490 ;
        RECT  10.400 3.900 10.640 4.620 ;
        RECT  7.870 4.380 10.640 4.620 ;
        RECT  14.630 1.580 14.870 3.780 ;
        RECT  14.550 3.380 16.260 3.780 ;
        RECT  13.880 1.060 15.430 1.300 ;
        RECT  15.190 1.060 15.430 2.620 ;
        RECT  15.190 2.380 16.650 2.620 ;
        RECT  13.880 1.060 14.130 3.600 ;
        RECT  16.500 1.850 17.130 2.090 ;
        RECT  18.660 2.380 19.330 2.620 ;
        RECT  16.890 1.850 17.130 3.100 ;
        RECT  15.500 2.860 17.130 3.100 ;
        RECT  16.660 2.860 16.900 4.120 ;
        RECT  18.660 2.380 18.900 4.120 ;
        RECT  16.660 3.880 18.900 4.120 ;
    END
END sdprb2

MACRO sdprb1
    CLASS CORE ;
    FOREIGN sdprb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.296  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.580 7.630 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.257  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.460 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.264  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.180 3.390 19.610 3.710 ;
        RECT  19.180 1.370 19.460 3.710 ;
        RECT  18.680 1.370 19.460 1.610 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.111  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.500 3.390 18.340 3.630 ;
        RECT  17.500 1.210 17.780 3.630 ;
        RECT  17.200 1.210 17.780 1.530 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.520 0.460 2.460 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.090  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.550 4.120 6.020 4.520 ;
        RECT  5.740 3.700 6.020 4.520 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.460 2.480 13.100 2.720 ;
        RECT  12.460 2.020 12.740 2.720 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.160 5.600 ;
        RECT  18.470 4.390 18.870 5.600 ;
        RECT  17.200 4.390 17.600 5.600 ;
        RECT  15.200 4.020 15.600 5.600 ;
        RECT  12.400 4.380 12.800 5.600 ;
        RECT  11.050 4.380 11.450 5.600 ;
        RECT  7.220 4.560 7.620 5.600 ;
        RECT  6.180 4.710 6.580 5.600 ;
        RECT  4.870 3.130 5.110 5.600 ;
        RECT  1.900 4.660 2.300 5.600 ;
        RECT  0.430 4.570 0.830 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.160 0.740 ;
        RECT  17.940 0.000 18.340 1.030 ;
        RECT  15.840 0.000 16.080 1.640 ;
        RECT  11.470 0.000 11.710 1.970 ;
        RECT  7.570 0.000 7.970 0.900 ;
        RECT  6.180 0.000 6.580 0.900 ;
        RECT  4.610 0.000 5.010 0.900 ;
        RECT  1.900 0.000 2.300 0.990 ;
        RECT  1.180 0.000 1.420 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.040 0.940 1.280 ;
        RECT  0.700 1.040 0.940 4.230 ;
        RECT  0.430 3.910 0.940 4.230 ;
        RECT  2.540 1.750 2.940 2.070 ;
        RECT  2.700 1.750 2.940 3.690 ;
        RECT  2.540 3.370 2.940 3.690 ;
        RECT  1.210 1.750 1.450 4.230 ;
        RECT  1.210 3.990 3.430 4.230 ;
        RECT  3.030 3.990 3.430 4.390 ;
        RECT  4.020 1.750 4.420 2.070 ;
        RECT  4.020 1.750 4.260 3.690 ;
        RECT  4.020 3.370 4.420 3.690 ;
        RECT  5.350 1.690 5.880 2.010 ;
        RECT  4.510 2.380 5.590 2.620 ;
        RECT  5.350 1.690 5.590 3.370 ;
        RECT  5.350 3.130 5.930 3.370 ;
        RECT  5.870 2.370 6.500 2.610 ;
        RECT  6.260 1.620 6.500 4.370 ;
        RECT  3.360 1.140 9.300 1.380 ;
        RECT  8.870 1.140 9.300 1.640 ;
        RECT  9.060 1.140 9.300 3.600 ;
        RECT  3.360 1.140 3.600 3.690 ;
        RECT  8.360 1.920 8.660 4.140 ;
        RECT  8.360 3.900 9.630 4.140 ;
        RECT  10.350 1.580 10.750 1.980 ;
        RECT  10.460 1.580 10.700 3.600 ;
        RECT  10.460 3.200 10.860 3.600 ;
        RECT  9.610 1.100 11.230 1.340 ;
        RECT  9.610 1.100 10.040 1.850 ;
        RECT  10.990 1.100 11.230 2.450 ;
        RECT  10.990 2.210 12.220 2.450 ;
        RECT  11.980 2.210 12.220 2.800 ;
        RECT  9.800 1.100 10.040 3.600 ;
        RECT  13.030 1.580 13.580 1.900 ;
        RECT  10.950 2.720 11.540 2.960 ;
        RECT  11.300 2.720 11.540 3.600 ;
        RECT  13.340 1.580 13.580 3.600 ;
        RECT  11.300 3.200 13.580 3.600 ;
        RECT  6.980 1.920 8.110 2.160 ;
        RECT  6.980 3.280 8.110 3.520 ;
        RECT  10.400 3.900 13.880 4.140 ;
        RECT  7.870 1.920 8.110 4.620 ;
        RECT  13.640 3.900 13.880 4.490 ;
        RECT  10.400 3.900 10.640 4.620 ;
        RECT  7.870 4.380 10.640 4.620 ;
        RECT  14.630 1.580 14.870 3.780 ;
        RECT  14.550 3.380 16.260 3.780 ;
        RECT  13.880 1.060 15.430 1.300 ;
        RECT  15.190 1.060 15.430 2.620 ;
        RECT  15.190 2.380 16.650 2.620 ;
        RECT  13.880 1.060 14.130 3.600 ;
        RECT  16.500 1.850 17.130 2.090 ;
        RECT  16.890 1.850 17.130 3.100 ;
        RECT  15.500 2.860 17.130 3.100 ;
        RECT  16.660 2.860 16.900 4.120 ;
        RECT  18.580 2.710 18.820 4.120 ;
        RECT  16.660 3.880 18.820 4.120 ;
    END
END sdprb1

MACRO sdpfb4
    CLASS CORE ;
    FOREIGN sdpfb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.010 2.520 5.530 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.453  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.120 2.830 ;
        RECT  3.880 2.150 4.120 2.830 ;
        RECT  3.420 2.580 3.860 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.014  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.980 3.150 15.290 3.390 ;
        RECT  14.930 1.450 15.170 2.030 ;
        RECT  13.250 1.830 15.170 2.030 ;
        RECT  13.450 1.790 15.170 2.030 ;
        RECT  13.450 1.420 13.690 2.130 ;
        RECT  12.940 2.020 13.470 2.460 ;
        RECT  12.980 2.020 13.220 3.390 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.897  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.850 2.930 19.600 3.170 ;
        RECT  17.850 1.680 19.570 1.920 ;
        RECT  19.330 1.310 19.570 1.920 ;
        RECT  17.850 2.550 18.250 3.250 ;
        RECT  17.850 1.150 18.090 3.250 ;
        RECT  17.420 2.020 18.090 2.460 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.240 2.550 0.640 2.950 ;
        RECT  0.240 2.020 0.500 2.950 ;
        RECT  0.120 2.020 0.500 2.460 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.020 1.590 3.560 1.990 ;
        RECT  2.000 2.130 3.260 2.370 ;
        RECT  3.020 1.590 3.260 2.370 ;
        RECT  2.240 3.140 2.740 3.580 ;
        RECT  2.500 2.130 2.740 3.580 ;
        RECT  2.000 2.130 2.240 2.710 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.140 2.020 10.640 2.620 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 22.960 5.600 ;
        RECT  19.790 4.590 20.190 5.600 ;
        RECT  18.430 4.590 18.830 5.600 ;
        RECT  16.890 4.590 17.290 5.600 ;
        RECT  15.480 4.630 15.880 5.600 ;
        RECT  14.120 4.630 14.520 5.600 ;
        RECT  12.550 4.600 12.960 5.600 ;
        RECT  11.020 4.160 11.420 5.600 ;
        RECT  9.620 4.260 10.020 5.600 ;
        RECT  7.800 4.770 8.210 5.600 ;
        RECT  6.090 4.420 6.510 5.600 ;
        RECT  4.820 4.390 5.220 5.600 ;
        RECT  2.280 4.380 2.680 5.600 ;
        RECT  0.910 4.380 1.310 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 22.960 0.740 ;
        RECT  19.990 0.000 20.390 1.440 ;
        RECT  18.510 0.000 18.910 1.440 ;
        RECT  17.030 0.000 17.430 1.450 ;
        RECT  15.590 0.000 15.990 1.550 ;
        RECT  14.110 0.000 14.510 1.550 ;
        RECT  12.620 0.000 13.030 1.650 ;
        RECT  9.460 0.000 9.860 1.200 ;
        RECT  5.590 0.000 5.990 0.890 ;
        RECT  4.660 0.000 5.060 0.890 ;
        RECT  2.230 0.000 2.640 1.230 ;
        RECT  0.930 0.000 1.330 0.900 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.460 1.240 1.700 ;
        RECT  1.000 1.460 1.240 4.040 ;
        RECT  0.150 3.800 1.240 4.040 ;
        RECT  1.480 1.490 1.920 1.890 ;
        RECT  1.480 1.650 2.780 1.890 ;
        RECT  1.480 1.490 1.720 3.120 ;
        RECT  1.560 2.940 1.800 3.520 ;
        RECT  6.500 2.290 7.340 2.530 ;
        RECT  6.500 1.630 6.740 3.450 ;
        RECT  6.500 3.210 7.250 3.450 ;
        RECT  6.550 0.980 7.560 1.220 ;
        RECT  3.430 1.110 4.010 1.350 ;
        RECT  3.870 1.130 6.790 1.370 ;
        RECT  7.320 0.980 7.560 2.040 ;
        RECT  7.320 1.800 8.020 2.040 ;
        RECT  7.780 1.800 8.020 3.400 ;
        RECT  3.500 3.730 4.610 3.970 ;
        RECT  4.370 1.130 4.610 3.980 ;
        RECT  5.040 1.610 6.260 1.850 ;
        RECT  5.040 1.610 5.280 2.170 ;
        RECT  6.020 1.610 6.260 4.060 ;
        RECT  5.530 3.820 7.350 4.060 ;
        RECT  7.110 3.820 7.350 4.420 ;
        RECT  7.110 4.180 8.220 4.420 ;
        RECT  8.800 1.120 9.040 1.640 ;
        RECT  8.750 1.460 8.990 2.980 ;
        RECT  8.750 2.740 9.350 2.980 ;
        RECT  9.110 2.740 9.350 3.400 ;
        RECT  7.950 1.130 8.510 1.530 ;
        RECT  8.260 1.130 8.510 3.900 ;
        RECT  8.260 3.500 8.680 3.900 ;
        RECT  9.630 3.490 11.300 3.730 ;
        RECT  11.060 2.280 11.300 3.730 ;
        RECT  8.260 3.660 9.870 3.900 ;
        RECT  15.370 2.180 16.610 2.580 ;
        RECT  16.370 1.410 16.610 3.270 ;
        RECT  10.810 0.980 12.330 1.220 ;
        RECT  10.810 0.980 11.050 1.720 ;
        RECT  9.640 1.480 11.050 1.720 ;
        RECT  20.770 1.010 21.010 1.790 ;
        RECT  9.230 2.150 9.880 2.390 ;
        RECT  12.090 0.980 12.330 3.230 ;
        RECT  9.640 1.480 9.880 3.250 ;
        RECT  12.090 2.990 12.700 3.230 ;
        RECT  9.640 3.010 10.800 3.250 ;
        RECT  12.460 2.990 12.700 3.870 ;
        RECT  20.650 1.550 20.890 3.870 ;
        RECT  12.460 3.630 20.890 3.870 ;
        RECT  21.250 1.050 21.830 1.290 ;
        RECT  21.250 1.050 21.490 1.960 ;
        RECT  21.420 1.720 21.660 4.130 ;
        RECT  11.510 1.570 11.750 2.110 ;
        RECT  11.540 1.970 11.780 3.720 ;
        RECT  11.540 3.480 12.110 3.720 ;
        RECT  22.100 1.750 22.340 3.760 ;
        RECT  11.870 3.480 12.110 4.350 ;
        RECT  11.870 4.110 20.890 4.350 ;
        RECT  20.650 4.110 20.890 4.620 ;
        RECT  22.160 3.520 22.400 4.620 ;
        RECT  20.650 4.380 22.400 4.620 ;
    END
END sdpfb4

MACRO sdpfb2
    CLASS CORE ;
    FOREIGN sdpfb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.010 2.520 5.530 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.453  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.120 2.830 ;
        RECT  3.880 2.150 4.120 2.830 ;
        RECT  3.420 2.580 3.860 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.614  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.980 3.150 13.740 3.390 ;
        RECT  13.450 1.420 13.690 2.090 ;
        RECT  12.940 2.020 13.520 2.460 ;
        RECT  13.250 1.830 13.690 2.090 ;
        RECT  12.980 2.020 13.220 3.390 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.511  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.460 2.550 16.700 3.250 ;
        RECT  16.380 1.150 16.620 2.750 ;
        RECT  15.740 2.020 16.620 2.460 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.240 2.550 0.640 2.950 ;
        RECT  0.240 2.020 0.500 2.950 ;
        RECT  0.120 2.020 0.500 2.460 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.478  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.020 1.590 3.560 1.910 ;
        RECT  2.000 2.130 3.260 2.370 ;
        RECT  3.020 1.590 3.260 2.370 ;
        RECT  2.240 3.140 2.740 3.580 ;
        RECT  2.500 2.130 2.740 3.580 ;
        RECT  2.000 2.130 2.240 2.710 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.140 2.020 10.640 2.620 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.160 5.600 ;
        RECT  16.960 4.590 17.360 5.600 ;
        RECT  15.420 4.590 15.820 5.600 ;
        RECT  14.120 4.630 14.520 5.600 ;
        RECT  12.550 4.600 12.960 5.600 ;
        RECT  11.020 4.160 11.420 5.600 ;
        RECT  9.620 4.260 10.020 5.600 ;
        RECT  7.800 4.770 8.210 5.600 ;
        RECT  6.090 4.420 6.510 5.600 ;
        RECT  4.820 4.390 5.220 5.600 ;
        RECT  2.280 4.380 2.680 5.600 ;
        RECT  0.910 4.380 1.310 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.160 0.740 ;
        RECT  17.040 0.000 17.440 1.440 ;
        RECT  15.560 0.000 15.960 1.450 ;
        RECT  14.110 0.000 14.510 1.550 ;
        RECT  12.620 0.000 13.030 1.650 ;
        RECT  9.460 0.000 9.860 1.200 ;
        RECT  5.590 0.000 5.990 0.890 ;
        RECT  4.660 0.000 5.060 0.890 ;
        RECT  2.230 0.000 2.640 1.230 ;
        RECT  0.930 0.000 1.330 0.900 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.460 1.240 1.700 ;
        RECT  1.000 1.460 1.240 4.040 ;
        RECT  0.150 3.800 1.240 4.040 ;
        RECT  1.480 1.490 1.920 1.890 ;
        RECT  1.480 1.650 2.780 1.890 ;
        RECT  1.480 1.490 1.720 3.120 ;
        RECT  1.560 2.940 1.800 3.520 ;
        RECT  6.500 2.290 7.340 2.530 ;
        RECT  6.500 1.630 6.740 3.450 ;
        RECT  6.500 3.210 7.250 3.450 ;
        RECT  6.550 0.980 7.560 1.220 ;
        RECT  3.430 1.110 4.010 1.350 ;
        RECT  3.870 1.130 6.790 1.370 ;
        RECT  7.320 0.980 7.560 2.040 ;
        RECT  7.320 1.800 8.020 2.040 ;
        RECT  7.780 1.800 8.020 3.400 ;
        RECT  4.370 1.130 4.610 3.750 ;
        RECT  3.310 3.510 4.610 3.750 ;
        RECT  5.040 1.610 6.260 1.850 ;
        RECT  5.040 1.610 5.280 2.170 ;
        RECT  6.020 1.610 6.260 4.060 ;
        RECT  5.530 3.820 7.350 4.060 ;
        RECT  7.110 3.820 7.350 4.420 ;
        RECT  7.110 4.180 8.220 4.420 ;
        RECT  8.800 1.120 9.040 1.640 ;
        RECT  8.750 1.460 8.990 2.980 ;
        RECT  8.750 2.740 9.350 2.980 ;
        RECT  9.110 2.740 9.350 3.400 ;
        RECT  7.950 1.130 8.510 1.530 ;
        RECT  8.260 1.130 8.510 3.900 ;
        RECT  8.260 3.500 8.680 3.900 ;
        RECT  9.630 3.490 11.300 3.730 ;
        RECT  11.060 2.280 11.300 3.730 ;
        RECT  8.260 3.660 9.870 3.900 ;
        RECT  13.900 2.240 15.140 2.640 ;
        RECT  14.900 1.410 15.140 3.390 ;
        RECT  10.810 0.980 12.330 1.220 ;
        RECT  10.810 0.980 11.050 1.720 ;
        RECT  9.640 1.480 11.050 1.720 ;
        RECT  17.850 1.010 18.090 1.790 ;
        RECT  9.230 2.150 9.880 2.390 ;
        RECT  12.090 0.980 12.330 3.230 ;
        RECT  9.640 1.480 9.880 3.250 ;
        RECT  12.090 2.990 12.700 3.230 ;
        RECT  9.640 3.010 10.800 3.250 ;
        RECT  12.460 2.990 12.700 3.870 ;
        RECT  17.730 1.550 17.970 3.870 ;
        RECT  12.460 3.630 17.970 3.870 ;
        RECT  18.330 1.050 18.910 1.290 ;
        RECT  18.330 1.050 18.570 1.960 ;
        RECT  18.500 1.720 18.740 4.130 ;
        RECT  11.510 1.570 11.750 2.110 ;
        RECT  11.540 1.970 11.780 3.720 ;
        RECT  11.540 3.480 12.110 3.720 ;
        RECT  19.180 1.750 19.420 3.760 ;
        RECT  11.870 3.480 12.110 4.350 ;
        RECT  11.870 4.110 17.970 4.350 ;
        RECT  17.730 4.110 17.970 4.620 ;
        RECT  19.240 3.520 19.480 4.620 ;
        RECT  17.730 4.380 19.480 4.620 ;
    END
END sdpfb2

MACRO sdpfb1
    CLASS CORE ;
    FOREIGN sdpfb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.520 5.530 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.660 2.210 4.340 2.450 ;
        RECT  3.940 1.990 4.340 2.450 ;
        RECT  3.420 2.580 3.920 3.020 ;
        RECT  3.660 2.210 3.920 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.067  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.320 1.890 13.330 2.130 ;
        RECT  13.090 1.420 13.330 2.130 ;
        RECT  12.320 3.010 13.100 3.250 ;
        RECT  12.320 1.890 12.820 2.460 ;
        RECT  12.320 1.890 12.620 3.250 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.294  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.090 1.070 15.600 1.470 ;
        RECT  14.620 2.930 15.330 3.170 ;
        RECT  14.620 2.020 15.330 2.460 ;
        RECT  15.090 1.070 15.330 2.460 ;
        RECT  14.620 2.020 14.860 3.170 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        RECT  1.990 2.450 2.740 2.690 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.530 2.020 10.020 2.620 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.920 5.600 ;
        RECT  14.060 4.380 14.300 5.600 ;
        RECT  11.920 4.600 12.320 5.600 ;
        RECT  10.360 4.340 10.780 5.600 ;
        RECT  8.970 4.260 9.380 5.600 ;
        RECT  7.070 4.770 7.470 5.600 ;
        RECT  5.500 4.420 5.900 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.720 3.550 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.920 0.740 ;
        RECT  14.450 0.000 14.850 1.450 ;
        RECT  12.270 0.000 12.670 1.650 ;
        RECT  9.340 0.000 9.740 1.200 ;
        RECT  5.590 0.000 5.990 0.890 ;
        RECT  3.270 0.000 3.670 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.250 1.750 ;
        RECT  1.010 1.510 1.250 3.310 ;
        RECT  0.230 3.070 1.250 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.510 1.570 1.910 2.210 ;
        RECT  1.510 1.970 3.420 2.210 ;
        RECT  1.510 1.570 1.750 4.440 ;
        RECT  1.510 3.950 1.800 4.440 ;
        RECT  6.420 1.610 6.820 2.030 ;
        RECT  6.580 2.210 7.130 2.610 ;
        RECT  6.580 1.610 6.820 3.210 ;
        RECT  6.320 2.970 6.820 3.210 ;
        RECT  6.320 2.970 6.560 3.530 ;
        RECT  5.080 1.660 5.320 2.280 ;
        RECT  5.080 2.040 6.080 2.280 ;
        RECT  5.840 2.320 6.340 2.720 ;
        RECT  5.840 2.040 6.080 4.060 ;
        RECT  4.920 3.820 6.820 4.060 ;
        RECT  6.580 3.820 6.820 4.530 ;
        RECT  6.580 4.290 7.600 4.530 ;
        RECT  4.460 0.980 4.870 1.370 ;
        RECT  2.070 0.980 2.770 1.220 ;
        RECT  6.550 0.980 7.520 1.220 ;
        RECT  4.460 1.130 6.790 1.370 ;
        RECT  2.530 0.980 2.770 1.730 ;
        RECT  7.120 0.980 7.520 1.600 ;
        RECT  4.460 0.980 4.820 1.730 ;
        RECT  2.530 1.490 4.820 1.730 ;
        RECT  4.580 0.980 4.820 2.940 ;
        RECT  7.370 1.380 7.610 3.330 ;
        RECT  7.060 2.930 7.610 3.330 ;
        RECT  4.320 2.690 4.610 3.670 ;
        RECT  4.210 3.210 4.610 3.670 ;
        RECT  1.990 3.430 4.610 3.670 ;
        RECT  8.500 0.980 9.000 1.330 ;
        RECT  8.500 0.980 8.940 1.380 ;
        RECT  8.500 0.980 8.740 1.930 ;
        RECT  8.330 1.690 8.570 3.410 ;
        RECT  8.330 3.000 8.790 3.410 ;
        RECT  7.850 1.010 8.260 1.420 ;
        RECT  10.410 2.440 10.650 3.970 ;
        RECT  7.630 3.730 10.650 3.970 ;
        RECT  7.850 1.010 8.090 4.040 ;
        RECT  7.630 3.630 8.090 4.040 ;
        RECT  13.220 2.370 14.030 2.620 ;
        RECT  13.790 1.410 14.030 3.170 ;
        RECT  13.400 2.930 14.030 3.170 ;
        RECT  10.290 0.980 11.940 1.220 ;
        RECT  9.120 1.540 10.530 1.780 ;
        RECT  10.290 0.980 10.530 1.780 ;
        RECT  15.970 1.010 16.210 1.950 ;
        RECT  15.570 1.710 16.210 1.950 ;
        RECT  9.050 1.610 9.290 3.270 ;
        RECT  8.810 2.280 9.290 2.690 ;
        RECT  9.040 2.280 9.290 3.270 ;
        RECT  9.040 3.030 10.150 3.270 ;
        RECT  11.700 0.980 11.940 3.730 ;
        RECT  13.290 3.420 15.810 3.660 ;
        RECT  11.700 3.490 13.480 3.730 ;
        RECT  15.570 1.710 15.810 4.130 ;
        RECT  16.460 1.050 17.030 1.290 ;
        RECT  16.460 1.050 16.700 2.450 ;
        RECT  16.050 2.210 16.710 2.450 ;
        RECT  16.050 2.210 16.300 4.050 ;
        RECT  16.050 3.810 16.670 4.050 ;
        RECT  11.150 1.650 11.390 3.530 ;
        RECT  17.440 1.750 17.700 3.580 ;
        RECT  17.090 3.340 17.700 3.580 ;
        RECT  11.220 2.130 11.460 4.350 ;
        RECT  12.360 3.970 15.020 4.140 ;
        RECT  13.660 3.900 15.020 4.140 ;
        RECT  11.220 4.110 13.850 4.220 ;
        RECT  11.220 4.110 12.760 4.350 ;
        RECT  14.720 3.900 15.020 4.620 ;
        RECT  17.090 3.340 17.330 4.620 ;
        RECT  14.720 4.380 17.330 4.620 ;
    END
END sdpfb1

MACRO sdnrq4
    CLASS CORE ;
    FOREIGN sdnrq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.110 2.340 15.560 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.660 2.210 4.340 2.450 ;
        RECT  3.940 1.990 4.340 2.450 ;
        RECT  3.420 2.580 3.920 3.020 ;
        RECT  3.660 2.210 3.920 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.006  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.130 1.440 12.060 1.680 ;
        RECT  11.660 1.060 12.060 1.680 ;
        RECT  9.870 2.970 11.650 3.210 ;
        RECT  9.870 2.880 10.580 3.290 ;
        RECT  10.130 1.440 10.580 3.290 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        RECT  1.990 2.450 2.740 2.690 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.680 5.600 ;
        RECT  14.560 4.300 14.960 5.600 ;
        RECT  12.020 4.710 12.420 5.600 ;
        RECT  10.660 4.710 11.060 5.600 ;
        RECT  9.120 4.710 9.520 5.600 ;
        RECT  6.290 4.240 6.690 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.800 3.550 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.680 0.740 ;
        RECT  14.390 0.000 14.790 1.620 ;
        RECT  13.130 0.000 13.530 1.120 ;
        RECT  10.920 0.000 11.320 1.200 ;
        RECT  9.440 0.000 9.840 1.200 ;
        RECT  7.370 0.000 7.770 0.910 ;
        RECT  3.270 0.000 3.670 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.250 1.750 ;
        RECT  1.010 1.510 1.250 3.310 ;
        RECT  0.230 3.070 1.250 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.510 1.570 1.910 2.210 ;
        RECT  1.510 1.970 3.420 2.210 ;
        RECT  1.510 1.570 1.750 3.840 ;
        RECT  1.280 3.600 1.520 4.600 ;
        RECT  1.280 4.360 1.860 4.600 ;
        RECT  1.980 0.980 2.770 1.220 ;
        RECT  2.530 0.980 2.770 1.730 ;
        RECT  4.530 1.040 4.820 1.730 ;
        RECT  2.530 1.490 4.820 1.730 ;
        RECT  4.580 1.040 4.820 2.940 ;
        RECT  4.320 2.690 4.610 3.670 ;
        RECT  4.210 3.210 4.610 3.670 ;
        RECT  1.990 3.430 4.610 3.670 ;
        RECT  5.540 1.560 6.380 1.800 ;
        RECT  5.540 1.560 5.780 2.930 ;
        RECT  5.770 2.690 6.010 3.510 ;
        RECT  5.060 1.080 7.030 1.320 ;
        RECT  6.790 1.080 7.030 2.940 ;
        RECT  5.060 1.080 5.300 3.580 ;
        RECT  4.950 3.170 5.350 3.580 ;
        RECT  7.350 1.310 7.740 1.710 ;
        RECT  6.020 2.040 6.500 2.450 ;
        RECT  6.260 2.040 6.500 3.510 ;
        RECT  7.350 1.310 7.590 3.510 ;
        RECT  6.260 3.180 7.590 3.510 ;
        RECT  8.780 0.990 9.020 2.910 ;
        RECT  8.840 2.670 9.080 3.500 ;
        RECT  8.500 3.230 9.080 3.500 ;
        RECT  11.890 1.970 12.680 2.210 ;
        RECT  12.440 1.450 12.680 2.210 ;
        RECT  11.240 2.170 12.210 2.590 ;
        RECT  11.890 1.970 12.210 3.260 ;
        RECT  11.890 3.020 13.190 3.260 ;
        RECT  12.570 2.450 13.670 2.690 ;
        RECT  8.190 1.730 8.430 2.990 ;
        RECT  7.830 2.750 8.430 2.990 ;
        RECT  7.830 2.750 8.090 3.980 ;
        RECT  13.430 2.450 13.670 3.980 ;
        RECT  7.830 3.740 13.670 3.980 ;
        RECT  13.650 1.480 14.150 1.880 ;
        RECT  5.540 3.750 7.530 3.990 ;
        RECT  7.290 3.750 7.530 4.470 ;
        RECT  13.910 1.480 14.150 4.470 ;
        RECT  7.290 4.230 14.150 4.470 ;
        RECT  5.540 3.750 5.780 4.620 ;
        RECT  4.740 4.380 5.780 4.620 ;
        RECT  15.210 1.260 15.450 2.100 ;
        RECT  14.390 1.860 15.450 2.100 ;
        RECT  14.390 1.860 14.640 3.520 ;
        RECT  14.390 3.260 15.530 3.520 ;
    END
END sdnrq4

MACRO sdnrq2
    CLASS CORE ;
    FOREIGN sdnrq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.296  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.580 7.630 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.257  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.460 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.237  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.110 3.130 16.660 3.450 ;
        RECT  16.380 1.490 16.660 3.450 ;
        RECT  16.240 1.490 16.660 1.810 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.520 0.460 2.460 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.090  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.550 4.120 6.020 4.520 ;
        RECT  5.740 3.700 6.020 4.520 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.360 5.600 ;
        RECT  16.670 4.160 17.070 5.600 ;
        RECT  15.340 4.420 15.740 5.600 ;
        RECT  14.190 4.090 14.430 5.600 ;
        RECT  11.310 4.380 11.550 5.600 ;
        RECT  7.220 4.560 7.620 5.600 ;
        RECT  6.180 4.710 6.580 5.600 ;
        RECT  4.870 3.130 5.110 5.600 ;
        RECT  1.900 4.660 2.300 5.600 ;
        RECT  0.430 4.570 0.830 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.360 0.740 ;
        RECT  16.800 0.000 17.200 1.110 ;
        RECT  15.500 0.000 15.900 1.110 ;
        RECT  14.200 0.000 14.600 0.890 ;
        RECT  11.470 0.000 11.710 1.890 ;
        RECT  7.570 0.000 7.970 0.900 ;
        RECT  6.180 0.000 6.580 0.900 ;
        RECT  4.610 0.000 5.010 0.900 ;
        RECT  1.900 0.000 2.300 0.990 ;
        RECT  1.180 0.000 1.420 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.040 0.940 1.280 ;
        RECT  0.700 1.040 0.940 4.230 ;
        RECT  0.430 3.910 0.940 4.230 ;
        RECT  2.540 1.750 2.940 2.070 ;
        RECT  2.700 1.750 2.940 3.690 ;
        RECT  2.540 3.370 2.940 3.690 ;
        RECT  1.210 1.750 1.450 4.230 ;
        RECT  1.210 3.990 3.430 4.230 ;
        RECT  3.030 3.990 3.430 4.390 ;
        RECT  4.020 1.750 4.420 2.070 ;
        RECT  4.020 1.750 4.260 3.690 ;
        RECT  4.020 3.370 4.420 3.690 ;
        RECT  5.350 1.690 5.880 2.010 ;
        RECT  4.510 2.380 5.590 2.620 ;
        RECT  5.350 1.690 5.590 3.370 ;
        RECT  5.350 3.130 5.930 3.370 ;
        RECT  5.870 2.370 6.500 2.610 ;
        RECT  6.260 1.620 6.500 4.370 ;
        RECT  3.360 1.140 9.360 1.380 ;
        RECT  8.870 1.140 9.360 1.560 ;
        RECT  9.060 1.140 9.360 3.600 ;
        RECT  3.360 1.140 3.600 3.690 ;
        RECT  6.980 1.920 8.110 2.160 ;
        RECT  6.980 3.280 8.110 3.520 ;
        RECT  7.870 1.920 8.110 4.620 ;
        RECT  7.870 4.380 10.370 4.620 ;
        RECT  10.350 1.580 10.750 1.980 ;
        RECT  10.460 1.580 10.700 3.600 ;
        RECT  10.460 3.280 10.860 3.600 ;
        RECT  9.610 1.100 11.230 1.340 ;
        RECT  9.610 1.100 10.040 1.770 ;
        RECT  10.990 1.100 11.230 2.450 ;
        RECT  10.990 2.210 12.020 2.450 ;
        RECT  9.800 1.100 10.040 3.600 ;
        RECT  12.130 1.580 12.530 1.900 ;
        RECT  10.950 2.720 12.530 2.960 ;
        RECT  12.260 1.580 12.530 2.990 ;
        RECT  12.080 2.720 12.320 3.600 ;
        RECT  8.360 1.920 8.660 4.140 ;
        RECT  8.360 3.900 13.310 4.140 ;
        RECT  13.070 3.900 13.310 4.490 ;
        RECT  13.430 1.660 14.010 1.900 ;
        RECT  13.430 1.660 13.670 3.670 ;
        RECT  13.430 3.350 13.920 3.670 ;
        RECT  12.950 1.070 13.740 1.310 ;
        RECT  13.500 1.180 14.490 1.420 ;
        RECT  14.250 1.180 14.490 2.430 ;
        RECT  14.250 2.190 15.120 2.430 ;
        RECT  12.950 1.070 13.190 3.600 ;
        RECT  12.740 3.280 13.190 3.600 ;
        RECT  14.970 1.660 15.600 1.900 ;
        RECT  15.360 2.100 16.080 2.340 ;
        RECT  15.360 1.660 15.600 2.910 ;
        RECT  14.010 2.670 15.600 2.910 ;
        RECT  14.890 2.670 15.130 3.450 ;
    END
END sdnrq2

MACRO sdnrq1
    CLASS CORE ;
    FOREIGN sdnrq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.296  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.580 7.630 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.257  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.460 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.189  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.110 3.130 16.660 3.450 ;
        RECT  16.380 1.490 16.660 3.450 ;
        RECT  16.240 1.490 16.660 1.810 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.520 0.460 2.460 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.090  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.550 4.120 6.020 4.520 ;
        RECT  5.740 3.700 6.020 4.520 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  15.500 4.420 15.900 5.600 ;
        RECT  14.190 4.090 14.430 5.600 ;
        RECT  11.310 4.380 11.550 5.600 ;
        RECT  7.220 4.560 7.620 5.600 ;
        RECT  6.180 4.710 6.580 5.600 ;
        RECT  4.870 3.130 5.110 5.600 ;
        RECT  1.900 4.660 2.300 5.600 ;
        RECT  0.430 4.570 0.830 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  15.500 0.000 15.900 1.110 ;
        RECT  14.200 0.000 14.600 0.890 ;
        RECT  11.470 0.000 11.710 1.890 ;
        RECT  7.570 0.000 7.970 0.900 ;
        RECT  6.180 0.000 6.580 0.900 ;
        RECT  4.610 0.000 5.010 0.900 ;
        RECT  1.900 0.000 2.300 0.990 ;
        RECT  1.180 0.000 1.420 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.040 0.940 1.280 ;
        RECT  0.700 1.040 0.940 4.230 ;
        RECT  0.430 3.910 0.940 4.230 ;
        RECT  2.540 1.750 2.940 2.070 ;
        RECT  2.700 1.750 2.940 3.690 ;
        RECT  2.540 3.370 2.940 3.690 ;
        RECT  1.210 1.750 1.450 4.230 ;
        RECT  1.210 3.990 3.430 4.230 ;
        RECT  3.030 3.990 3.430 4.390 ;
        RECT  4.020 1.750 4.420 2.070 ;
        RECT  4.020 1.750 4.260 3.690 ;
        RECT  4.020 3.370 4.420 3.690 ;
        RECT  5.350 1.690 5.880 2.010 ;
        RECT  4.510 2.380 5.590 2.620 ;
        RECT  5.350 1.690 5.590 3.370 ;
        RECT  5.350 3.130 5.930 3.370 ;
        RECT  5.870 2.370 6.500 2.610 ;
        RECT  6.260 1.620 6.500 4.370 ;
        RECT  3.360 1.140 9.360 1.380 ;
        RECT  8.870 1.140 9.360 1.560 ;
        RECT  9.060 1.140 9.360 3.600 ;
        RECT  3.360 1.140 3.600 3.690 ;
        RECT  6.980 1.920 8.110 2.160 ;
        RECT  6.980 3.280 8.110 3.520 ;
        RECT  7.870 1.920 8.110 4.620 ;
        RECT  7.870 4.380 10.370 4.620 ;
        RECT  10.350 1.580 10.750 1.980 ;
        RECT  10.460 1.580 10.700 3.600 ;
        RECT  10.460 3.280 10.860 3.600 ;
        RECT  9.610 1.100 11.230 1.340 ;
        RECT  9.610 1.100 10.040 1.770 ;
        RECT  10.990 1.100 11.230 2.450 ;
        RECT  10.990 2.210 12.020 2.450 ;
        RECT  9.800 1.100 10.040 3.600 ;
        RECT  12.130 1.580 12.500 1.900 ;
        RECT  10.950 2.720 12.500 2.960 ;
        RECT  12.260 1.580 12.500 2.990 ;
        RECT  12.080 2.720 12.320 3.600 ;
        RECT  8.360 1.920 8.660 4.140 ;
        RECT  8.360 3.900 13.310 4.140 ;
        RECT  13.070 3.900 13.310 4.490 ;
        RECT  13.430 1.660 14.010 1.900 ;
        RECT  13.430 1.660 13.670 3.670 ;
        RECT  13.430 3.350 13.920 3.670 ;
        RECT  12.950 1.070 13.840 1.310 ;
        RECT  13.600 1.180 14.490 1.420 ;
        RECT  14.250 1.180 14.490 2.430 ;
        RECT  14.250 2.190 15.120 2.430 ;
        RECT  12.950 1.070 13.190 3.600 ;
        RECT  12.740 3.280 13.190 3.600 ;
        RECT  14.970 1.660 15.600 1.900 ;
        RECT  15.360 2.100 16.080 2.340 ;
        RECT  15.360 1.660 15.600 2.910 ;
        RECT  14.010 2.670 15.600 2.910 ;
        RECT  14.890 2.670 15.130 3.450 ;
    END
END sdnrq1

MACRO sdnrn4
    CLASS CORE ;
    FOREIGN sdnrn4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.180 2.580 15.560 3.020 ;
        RECT  15.180 2.160 15.420 3.020 ;
        RECT  14.940 2.160 15.420 2.560 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.970 2.580 4.420 3.020 ;
        RECT  3.970 2.130 4.370 3.020 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.802  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.940 3.140 13.380 3.580 ;
        RECT  11.250 2.900 13.360 3.140 ;
        RECT  13.120 1.820 13.360 3.580 ;
        RECT  11.000 1.820 13.360 2.060 ;
        RECT  12.300 1.490 12.540 2.060 ;
        RECT  11.000 1.510 11.240 2.060 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.780 2.930 ;
        RECT  0.120 2.520 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.210 1.990 2.740 2.460 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.680 5.600 ;
        RECT  14.390 4.300 14.790 5.600 ;
        RECT  13.110 4.370 13.510 5.600 ;
        RECT  11.810 4.370 12.210 5.600 ;
        RECT  10.510 4.400 10.910 5.600 ;
        RECT  9.180 4.710 9.580 5.600 ;
        RECT  6.390 4.580 6.830 5.600 ;
        RECT  3.190 4.200 3.590 5.600 ;
        RECT  0.720 4.470 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.680 0.740 ;
        RECT  14.330 0.000 14.730 1.440 ;
        RECT  13.040 0.000 13.440 0.980 ;
        RECT  11.570 0.000 11.970 1.200 ;
        RECT  9.480 0.000 9.880 1.270 ;
        RECT  7.420 0.000 7.820 0.910 ;
        RECT  3.250 0.980 3.800 1.220 ;
        RECT  3.560 0.000 3.800 1.220 ;
        RECT  0.920 0.000 1.320 0.930 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.440 1.260 1.680 ;
        RECT  1.020 1.440 1.260 3.500 ;
        RECT  1.020 2.240 1.470 2.640 ;
        RECT  1.020 2.240 1.270 3.500 ;
        RECT  0.150 3.260 1.270 3.500 ;
        RECT  1.510 1.600 1.960 2.000 ;
        RECT  1.720 2.760 3.240 3.000 ;
        RECT  3.000 2.010 3.240 3.000 ;
        RECT  1.720 1.600 1.960 3.130 ;
        RECT  1.540 2.890 1.780 4.620 ;
        RECT  2.050 0.980 2.600 1.220 ;
        RECT  2.360 0.980 2.600 1.700 ;
        RECT  4.530 1.000 4.770 1.700 ;
        RECT  2.360 1.460 4.770 1.700 ;
        RECT  3.480 1.460 3.720 3.610 ;
        RECT  2.070 3.370 4.710 3.610 ;
        RECT  2.070 3.370 2.310 3.920 ;
        RECT  4.470 3.370 4.710 4.100 ;
        RECT  5.520 1.540 6.360 1.780 ;
        RECT  5.520 1.540 5.760 3.430 ;
        RECT  5.520 3.190 6.100 3.430 ;
        RECT  5.040 1.060 7.120 1.300 ;
        RECT  6.880 1.060 7.120 2.940 ;
        RECT  5.040 1.060 5.280 3.270 ;
        RECT  6.120 2.060 6.580 2.460 ;
        RECT  6.340 2.060 6.580 3.450 ;
        RECT  7.400 1.630 7.640 3.450 ;
        RECT  6.340 3.210 7.640 3.450 ;
        RECT  8.700 0.980 9.140 1.300 ;
        RECT  8.700 0.980 8.940 3.460 ;
        RECT  8.540 3.140 8.940 3.460 ;
        RECT  10.300 1.280 10.540 1.820 ;
        RECT  9.180 1.580 10.540 1.820 ;
        RECT  9.180 1.580 9.420 3.140 ;
        RECT  9.180 2.900 10.380 3.140 ;
        RECT  8.220 1.720 8.460 2.270 ;
        RECT  7.880 2.030 8.460 2.270 ;
        RECT  9.780 2.360 12.880 2.600 ;
        RECT  10.640 2.360 10.880 3.640 ;
        RECT  9.180 3.400 10.880 3.640 ;
        RECT  7.880 2.030 8.120 3.990 ;
        RECT  9.180 3.400 9.420 3.990 ;
        RECT  7.880 3.750 9.420 3.990 ;
        RECT  13.670 3.130 14.220 3.370 ;
        RECT  13.670 1.270 13.910 4.120 ;
        RECT  9.660 3.880 13.910 4.120 ;
        RECT  5.090 3.940 7.520 4.180 ;
        RECT  7.280 3.940 7.520 4.470 ;
        RECT  9.660 3.880 9.900 4.470 ;
        RECT  7.280 4.230 9.900 4.470 ;
        RECT  5.090 3.940 5.330 4.620 ;
        RECT  4.770 4.380 5.330 4.620 ;
        RECT  15.150 1.270 15.390 1.920 ;
        RECT  14.160 1.680 15.390 1.920 ;
        RECT  14.160 1.680 14.400 2.890 ;
        RECT  14.160 2.650 14.700 2.890 ;
        RECT  14.460 2.650 14.700 3.510 ;
        RECT  14.460 3.270 15.530 3.510 ;
    END
END sdnrn4

MACRO sdnrn2
    CLASS CORE ;
    FOREIGN sdnrn2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.415  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.220 1.460 16.740 1.900 ;
        RECT  16.220 1.460 16.470 3.450 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.360 5.600 ;
        RECT  16.890 4.170 17.130 5.600 ;
        RECT  15.590 4.170 15.830 5.600 ;
        RECT  14.310 3.990 14.550 5.600 ;
        RECT  11.290 4.350 11.530 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.360 0.740 ;
        RECT  16.810 0.000 17.210 1.010 ;
        RECT  15.510 0.000 15.910 1.010 ;
        RECT  14.020 0.000 14.420 0.890 ;
        RECT  11.280 0.000 11.520 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.560 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.150 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.150 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.510 4.110 ;
        RECT  10.320 1.750 10.560 3.610 ;
        RECT  10.320 3.290 10.740 3.610 ;
        RECT  9.580 1.270 11.040 1.510 ;
        RECT  10.800 1.270 11.040 2.600 ;
        RECT  10.800 2.360 12.040 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  11.940 1.830 12.520 2.070 ;
        RECT  12.280 1.830 12.520 3.100 ;
        RECT  10.940 2.860 12.520 3.100 ;
        RECT  11.810 2.860 12.050 3.630 ;
        RECT  11.810 3.390 12.380 3.630 ;
        RECT  9.850 3.870 12.010 4.110 ;
        RECT  11.770 3.870 12.010 4.580 ;
        RECT  11.770 4.340 12.740 4.580 ;
        RECT  13.450 1.610 13.840 1.930 ;
        RECT  13.450 1.610 13.690 4.040 ;
        RECT  13.450 3.720 13.860 4.040 ;
        RECT  12.760 1.130 14.590 1.370 ;
        RECT  14.350 1.130 14.590 2.530 ;
        RECT  14.560 2.290 14.960 2.690 ;
        RECT  12.760 1.130 13.000 3.180 ;
        RECT  12.800 2.940 13.040 3.710 ;
        RECT  14.830 1.780 15.440 2.020 ;
        RECT  13.940 2.770 14.180 3.390 ;
        RECT  15.200 1.780 15.440 3.390 ;
        RECT  13.940 3.150 15.440 3.390 ;
        RECT  14.890 3.150 15.130 3.720 ;
    END
END sdnrn2

MACRO sdnrn1
    CLASS CORE ;
    FOREIGN sdnrn1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.320 1.570 16.570 3.450 ;
        RECT  15.740 2.020 16.570 2.460 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  15.740 4.070 15.980 5.600 ;
        RECT  14.280 3.630 14.520 5.600 ;
        RECT  11.290 4.350 11.530 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  15.690 0.000 15.930 1.290 ;
        RECT  14.020 0.000 14.420 0.890 ;
        RECT  11.280 0.000 11.520 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.560 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.930 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.150 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.150 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.510 4.110 ;
        RECT  10.320 1.750 10.560 3.610 ;
        RECT  10.320 3.290 10.740 3.610 ;
        RECT  9.580 1.270 11.040 1.510 ;
        RECT  10.800 1.270 11.040 2.600 ;
        RECT  10.800 2.360 12.040 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  11.940 1.830 12.520 2.070 ;
        RECT  12.280 1.830 12.520 3.100 ;
        RECT  10.940 2.860 12.520 3.100 ;
        RECT  11.810 2.860 12.050 3.630 ;
        RECT  11.810 3.390 12.380 3.630 ;
        RECT  9.850 3.870 12.010 4.110 ;
        RECT  11.770 3.870 12.010 4.580 ;
        RECT  11.770 4.340 12.740 4.580 ;
        RECT  13.450 1.610 13.840 1.930 ;
        RECT  13.450 1.610 13.690 4.040 ;
        RECT  13.450 3.720 13.860 4.040 ;
        RECT  12.760 1.130 14.590 1.370 ;
        RECT  14.350 1.130 14.590 2.530 ;
        RECT  14.560 2.290 14.960 2.690 ;
        RECT  12.760 1.130 13.000 3.180 ;
        RECT  12.800 2.940 13.040 3.710 ;
        RECT  14.830 1.780 15.440 2.020 ;
        RECT  13.940 2.770 14.180 3.390 ;
        RECT  15.200 1.780 15.440 3.390 ;
        RECT  13.940 3.150 15.440 3.390 ;
        RECT  15.020 3.150 15.260 3.720 ;
    END
END sdnrn1

MACRO sdnrb4
    CLASS CORE ;
    FOREIGN sdnrb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.442  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.870 2.180 18.360 3.020 ;
        RECT  17.600 2.180 18.360 2.610 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.453  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.820 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.939  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.120 1.440 16.000 1.680 ;
        RECT  15.180 1.440 15.620 3.280 ;
        RECT  14.120 1.360 14.520 1.680 ;
        RECT  13.880 2.810 14.430 3.050 ;
        RECT  14.190 1.360 14.430 3.050 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.939  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.150 1.440 13.040 1.680 ;
        RECT  11.260 2.810 12.970 3.050 ;
        RECT  11.820 2.800 12.970 3.050 ;
        RECT  11.820 1.440 12.260 3.050 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.670 0.670 3.070 ;
        RECT  0.120 2.580 0.500 3.070 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.210 3.020 ;
        RECT  3.970 2.210 4.210 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 18.480 5.600 ;
        RECT  17.200 4.300 17.600 5.600 ;
        RECT  15.930 4.400 16.330 5.600 ;
        RECT  14.620 4.250 15.020 5.600 ;
        RECT  13.310 4.250 13.710 5.600 ;
        RECT  12.000 4.250 12.400 5.600 ;
        RECT  10.690 4.400 11.090 5.600 ;
        RECT  9.290 4.710 9.690 5.600 ;
        RECT  6.470 4.240 6.870 5.600 ;
        RECT  3.260 4.520 3.660 5.600 ;
        RECT  0.780 4.620 1.180 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 18.480 0.740 ;
        RECT  17.040 0.000 17.440 1.440 ;
        RECT  14.860 0.000 15.260 1.200 ;
        RECT  13.380 0.000 13.780 1.200 ;
        RECT  11.900 0.000 12.300 1.200 ;
        RECT  9.690 0.000 10.090 1.270 ;
        RECT  7.490 0.000 7.890 0.910 ;
        RECT  3.010 1.080 3.580 1.320 ;
        RECT  3.010 0.000 3.250 1.320 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.340 1.820 ;
        RECT  1.100 1.580 1.340 2.910 ;
        RECT  1.000 2.700 1.240 3.590 ;
        RECT  0.150 3.350 1.240 3.590 ;
        RECT  1.590 2.100 3.510 2.340 ;
        RECT  1.590 1.760 1.830 3.230 ;
        RECT  1.530 3.070 1.770 3.670 ;
        RECT  1.980 0.980 2.570 1.220 ;
        RECT  2.330 0.980 2.570 1.860 ;
        RECT  2.330 1.620 4.700 1.860 ;
        RECT  4.460 1.150 4.700 3.570 ;
        RECT  4.140 3.260 4.790 3.570 ;
        RECT  4.460 3.170 4.790 3.570 ;
        RECT  2.150 3.330 4.790 3.570 ;
        RECT  5.950 1.510 6.210 3.510 ;
        RECT  7.310 1.630 7.780 2.010 ;
        RECT  6.450 1.770 7.780 2.010 ;
        RECT  6.450 1.770 6.690 3.420 ;
        RECT  6.450 3.180 7.610 3.420 ;
        RECT  5.200 0.980 6.780 1.220 ;
        RECT  6.530 1.150 8.260 1.390 ;
        RECT  8.020 1.150 8.260 2.500 ;
        RECT  7.070 2.260 8.260 2.500 ;
        RECT  7.070 2.260 7.490 2.610 ;
        RECT  5.200 0.980 5.450 3.460 ;
        RECT  8.850 0.990 9.240 1.390 ;
        RECT  9.000 0.990 9.240 3.500 ;
        RECT  8.660 3.230 9.240 3.500 ;
        RECT  9.480 2.530 10.070 2.780 ;
        RECT  8.500 1.730 8.740 2.990 ;
        RECT  8.030 2.750 8.740 2.990 ;
        RECT  8.030 2.750 8.270 3.980 ;
        RECT  9.480 2.530 9.720 3.980 ;
        RECT  8.030 3.740 9.720 3.980 ;
        RECT  10.430 1.210 10.830 1.750 ;
        RECT  9.480 1.510 10.550 1.820 ;
        RECT  9.480 1.510 9.720 2.150 ;
        RECT  10.310 1.510 10.550 3.530 ;
        RECT  9.960 3.140 10.550 3.530 ;
        RECT  14.670 2.100 14.910 3.530 ;
        RECT  9.960 3.290 14.910 3.530 ;
        RECT  16.380 1.020 16.620 1.630 ;
        RECT  16.300 1.390 16.540 4.010 ;
        RECT  5.450 3.750 7.530 3.990 ;
        RECT  9.960 3.770 16.860 4.010 ;
        RECT  7.290 3.750 7.530 4.470 ;
        RECT  9.960 3.770 10.200 4.470 ;
        RECT  7.290 4.230 10.200 4.470 ;
        RECT  5.450 3.750 5.690 4.620 ;
        RECT  4.890 4.380 5.690 4.620 ;
        RECT  17.860 1.270 18.100 1.940 ;
        RECT  16.860 1.700 18.100 1.940 ;
        RECT  16.860 1.700 17.100 3.110 ;
        RECT  16.860 2.870 17.620 3.110 ;
        RECT  17.380 2.870 17.620 3.770 ;
        RECT  17.380 3.510 18.180 3.770 ;
    END
END sdnrb4

MACRO sdnrb2
    CLASS CORE ;
    FOREIGN sdnrb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.980 3.140 18.420 3.580 ;
        RECT  17.680 3.130 18.360 3.370 ;
        RECT  18.120 1.650 18.360 3.580 ;
        RECT  17.760 1.650 18.360 1.890 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.300 1.460 16.740 1.900 ;
        RECT  16.300 1.460 16.540 3.450 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.040 5.600 ;
        RECT  18.390 4.170 18.630 5.600 ;
        RECT  16.970 4.170 17.210 5.600 ;
        RECT  15.660 4.170 15.900 5.600 ;
        RECT  14.380 3.990 14.620 5.600 ;
        RECT  11.360 4.350 11.600 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.040 0.740 ;
        RECT  18.430 0.000 18.830 1.010 ;
        RECT  17.010 0.000 17.410 1.010 ;
        RECT  15.630 0.000 16.030 1.010 ;
        RECT  14.020 0.000 14.420 0.890 ;
        RECT  11.280 0.000 11.520 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.550 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.150 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.150 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.510 4.110 ;
        RECT  10.320 1.750 10.560 3.610 ;
        RECT  10.320 3.290 10.740 3.610 ;
        RECT  9.580 1.270 11.040 1.510 ;
        RECT  10.800 1.270 11.040 2.600 ;
        RECT  10.800 2.360 12.040 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  11.940 1.830 12.520 2.070 ;
        RECT  12.280 1.830 12.520 3.100 ;
        RECT  10.940 2.860 12.520 3.100 ;
        RECT  11.880 2.860 12.120 3.630 ;
        RECT  11.880 3.390 12.450 3.630 ;
        RECT  9.850 3.870 12.080 4.110 ;
        RECT  11.840 3.870 12.080 4.580 ;
        RECT  11.840 4.340 12.810 4.580 ;
        RECT  13.520 1.610 13.760 4.040 ;
        RECT  13.520 3.720 13.930 4.040 ;
        RECT  12.760 1.130 14.610 1.370 ;
        RECT  14.370 1.130 14.610 2.530 ;
        RECT  14.370 2.290 15.030 2.530 ;
        RECT  14.630 2.290 15.030 2.690 ;
        RECT  12.760 1.130 13.000 3.180 ;
        RECT  12.870 2.940 13.110 3.710 ;
        RECT  14.870 1.780 15.510 2.020 ;
        RECT  16.900 2.180 17.830 2.420 ;
        RECT  14.010 2.770 14.250 3.480 ;
        RECT  15.270 1.780 15.510 3.930 ;
        RECT  14.010 3.240 15.510 3.480 ;
        RECT  14.880 3.240 15.510 3.720 ;
        RECT  16.900 2.180 17.140 3.930 ;
        RECT  15.270 3.690 17.140 3.930 ;
    END
END sdnrb2

MACRO sdnrb1
    CLASS CORE ;
    FOREIGN sdnrb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.241  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.510 3.270 16.180 3.580 ;
        RECT  15.930 1.820 16.180 3.580 ;
        RECT  15.740 3.140 16.180 3.580 ;
        RECT  15.590 1.820 16.180 2.060 ;
        RECT  15.590 1.500 15.830 2.060 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.860 1.460 17.240 1.970 ;
        RECT  16.890 1.460 17.130 3.450 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.360 5.600 ;
        RECT  16.180 4.170 16.420 5.600 ;
        RECT  14.310 3.990 14.550 5.600 ;
        RECT  11.290 4.350 11.530 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.360 0.740 ;
        RECT  16.220 0.000 16.460 1.200 ;
        RECT  14.020 0.000 14.420 0.890 ;
        RECT  11.280 0.000 11.520 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.550 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.060 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.060 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.510 4.110 ;
        RECT  10.320 1.750 10.560 3.610 ;
        RECT  10.320 3.290 10.740 3.610 ;
        RECT  9.580 1.270 11.040 1.510 ;
        RECT  10.800 1.270 11.040 2.600 ;
        RECT  10.800 2.360 12.040 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  11.940 1.830 12.520 2.070 ;
        RECT  12.280 1.830 12.520 3.100 ;
        RECT  10.940 2.860 12.520 3.100 ;
        RECT  11.810 2.860 12.050 3.630 ;
        RECT  11.810 3.390 12.380 3.630 ;
        RECT  9.850 3.870 12.010 4.110 ;
        RECT  11.770 3.870 12.010 4.580 ;
        RECT  11.770 4.340 12.740 4.580 ;
        RECT  13.300 1.720 13.840 2.040 ;
        RECT  13.300 1.720 13.540 3.960 ;
        RECT  13.300 3.720 13.860 3.960 ;
        RECT  12.760 1.130 14.520 1.370 ;
        RECT  14.280 1.130 14.520 2.600 ;
        RECT  14.280 2.360 14.860 2.600 ;
        RECT  12.760 1.130 13.000 3.180 ;
        RECT  12.800 2.940 13.040 3.710 ;
        RECT  14.810 1.700 15.340 2.020 ;
        RECT  15.100 2.310 15.540 2.710 ;
        RECT  15.100 1.700 15.340 3.060 ;
        RECT  13.860 2.770 14.100 3.480 ;
        RECT  14.970 2.820 15.210 3.720 ;
        RECT  13.860 3.240 15.210 3.480 ;
        RECT  14.810 3.240 15.210 3.720 ;
    END
END sdnrb1

MACRO sdnfb4
    CLASS CORE ;
    FOREIGN sdnfb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.451  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.210 2.230 5.610 2.630 ;
        RECT  5.100 2.020 5.540 2.460 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.020 4.520 2.460 ;
        RECT  4.120 1.890 4.520 2.460 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.143  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.290 1.620 16.050 1.860 ;
        RECT  14.190 3.650 15.970 3.890 ;
        RECT  14.620 2.580 15.060 3.020 ;
        RECT  14.620 1.620 14.860 3.890 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.558  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.530 2.580 18.980 3.020 ;
        RECT  16.880 3.900 18.770 4.300 ;
        RECT  18.530 1.540 18.770 4.300 ;
        RECT  17.010 1.540 18.770 1.940 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.390 2.520 0.790 2.920 ;
        RECT  0.120 2.580 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.290 2.450 2.740 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.600 5.600 ;
        RECT  18.930 4.610 19.330 5.600 ;
        RECT  17.620 4.610 18.020 5.600 ;
        RECT  16.310 4.610 16.710 5.600 ;
        RECT  14.930 4.610 15.330 5.600 ;
        RECT  13.550 4.610 13.950 5.600 ;
        RECT  12.180 4.610 12.580 5.600 ;
        RECT  9.380 3.960 9.620 5.600 ;
        RECT  5.730 4.180 5.970 5.600 ;
        RECT  3.180 4.360 3.580 5.600 ;
        RECT  0.800 4.570 1.200 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.600 0.740 ;
        RECT  19.050 0.000 19.450 0.890 ;
        RECT  17.690 0.000 18.090 0.890 ;
        RECT  16.330 0.000 16.730 0.890 ;
        RECT  14.970 0.000 15.370 0.890 ;
        RECT  13.700 0.000 14.100 0.890 ;
        RECT  12.240 0.000 12.640 0.890 ;
        RECT  9.380 0.000 9.630 1.440 ;
        RECT  6.610 0.000 7.010 0.890 ;
        RECT  3.260 0.000 3.500 1.200 ;
        RECT  0.740 0.000 1.140 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.270 2.090 ;
        RECT  1.030 2.560 1.480 2.960 ;
        RECT  1.030 1.850 1.270 3.530 ;
        RECT  0.150 3.290 1.270 3.530 ;
        RECT  1.510 1.770 1.910 2.170 ;
        RECT  1.510 1.930 3.590 2.170 ;
        RECT  3.190 1.930 3.590 2.370 ;
        RECT  1.720 1.930 1.960 3.440 ;
        RECT  1.530 3.200 1.770 3.750 ;
        RECT  5.020 1.540 6.090 1.780 ;
        RECT  5.850 2.230 6.410 2.630 ;
        RECT  5.850 1.540 6.090 3.320 ;
        RECT  5.080 3.080 6.090 3.320 ;
        RECT  6.380 1.660 6.930 1.900 ;
        RECT  6.690 1.660 6.930 2.370 ;
        RECT  6.770 2.170 7.010 3.230 ;
        RECT  6.380 2.990 7.010 3.230 ;
        RECT  1.980 0.980 3.020 1.220 ;
        RECT  3.760 0.980 4.920 1.220 ;
        RECT  4.700 1.060 6.440 1.300 ;
        RECT  6.260 1.130 7.410 1.370 ;
        RECT  2.780 0.980 3.020 1.680 ;
        RECT  3.760 0.980 4.000 1.680 ;
        RECT  2.780 1.440 4.000 1.680 ;
        RECT  7.170 1.130 7.410 1.970 ;
        RECT  2.230 3.260 2.470 3.810 ;
        RECT  7.400 1.730 7.640 3.810 ;
        RECT  2.230 3.570 7.640 3.810 ;
        RECT  8.640 1.440 8.890 3.230 ;
        RECT  9.810 2.190 10.050 2.870 ;
        RECT  9.560 2.630 10.050 2.870 ;
        RECT  7.900 1.440 8.150 3.720 ;
        RECT  9.560 2.630 9.800 3.720 ;
        RECT  7.900 3.480 9.800 3.720 ;
        RECT  10.040 1.440 10.590 1.920 ;
        RECT  9.130 1.680 10.590 1.920 ;
        RECT  9.130 1.680 9.370 2.480 ;
        RECT  10.350 1.440 10.590 3.370 ;
        RECT  10.040 3.130 10.590 3.370 ;
        RECT  11.370 1.520 11.940 1.760 ;
        RECT  11.370 1.520 11.610 3.370 ;
        RECT  11.370 3.130 11.920 3.370 ;
        RECT  12.910 1.640 13.310 2.050 ;
        RECT  12.370 1.720 13.310 2.050 ;
        RECT  12.370 1.720 12.610 2.300 ;
        RECT  11.880 2.060 12.610 2.300 ;
        RECT  11.880 2.060 12.120 2.640 ;
        RECT  13.070 2.490 14.380 2.730 ;
        RECT  13.070 1.640 13.310 3.580 ;
        RECT  12.930 3.340 13.170 3.890 ;
        RECT  16.260 2.410 18.110 2.810 ;
        RECT  12.560 2.600 12.800 3.130 ;
        RECT  10.860 1.440 11.110 3.930 ;
        RECT  10.860 3.690 12.690 3.930 ;
        RECT  12.450 2.910 12.690 4.370 ;
        RECT  16.260 2.410 16.500 4.370 ;
        RECT  12.450 4.130 16.500 4.370 ;
    END
END sdnfb4

MACRO sdnfb2
    CLASS CORE ;
    FOREIGN sdnfb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.451  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.210 2.230 5.610 2.630 ;
        RECT  5.100 2.020 5.540 2.460 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.020 4.520 2.460 ;
        RECT  4.120 1.890 4.520 2.460 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.561  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.040 1.600 14.690 1.840 ;
        RECT  14.040 3.650 14.590 3.890 ;
        RECT  14.040 2.580 14.500 3.020 ;
        RECT  14.040 1.600 14.380 3.020 ;
        RECT  14.040 1.600 14.280 3.890 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.282  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.500 3.850 16.670 4.250 ;
        RECT  16.300 1.520 16.670 4.250 ;
        RECT  15.650 1.520 16.670 1.920 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.390 2.520 0.790 2.920 ;
        RECT  0.130 2.580 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.290 2.450 2.740 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  16.240 4.610 16.640 5.600 ;
        RECT  14.930 4.610 15.330 5.600 ;
        RECT  13.550 4.610 13.950 5.600 ;
        RECT  12.180 4.610 12.580 5.600 ;
        RECT  9.380 3.960 9.620 5.600 ;
        RECT  5.730 4.180 5.970 5.600 ;
        RECT  3.260 4.360 3.500 5.600 ;
        RECT  0.800 4.570 1.200 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  16.250 0.000 16.650 0.890 ;
        RECT  14.970 0.000 15.370 0.890 ;
        RECT  13.700 0.000 14.100 0.890 ;
        RECT  12.240 0.000 12.640 0.890 ;
        RECT  9.310 0.000 9.710 1.440 ;
        RECT  6.610 0.000 7.010 0.890 ;
        RECT  3.260 0.000 3.500 1.200 ;
        RECT  0.820 0.000 1.060 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.270 2.090 ;
        RECT  1.030 2.560 1.480 2.960 ;
        RECT  1.030 1.850 1.270 3.530 ;
        RECT  0.150 3.290 1.270 3.530 ;
        RECT  1.510 1.770 1.920 2.170 ;
        RECT  1.510 1.930 3.590 2.170 ;
        RECT  3.190 1.930 3.590 2.370 ;
        RECT  1.720 1.930 1.960 3.440 ;
        RECT  1.530 3.200 1.770 3.750 ;
        RECT  5.020 1.540 6.090 1.780 ;
        RECT  5.850 2.230 6.410 2.630 ;
        RECT  5.850 1.540 6.090 3.320 ;
        RECT  5.080 3.080 6.090 3.320 ;
        RECT  6.380 1.660 6.930 1.900 ;
        RECT  6.690 1.660 6.930 2.370 ;
        RECT  6.770 2.180 7.010 3.230 ;
        RECT  6.380 2.990 7.010 3.230 ;
        RECT  1.980 0.980 3.020 1.220 ;
        RECT  3.760 0.980 5.070 1.220 ;
        RECT  4.870 1.060 6.440 1.300 ;
        RECT  6.270 1.130 7.410 1.370 ;
        RECT  2.780 0.980 3.020 1.680 ;
        RECT  3.760 0.980 4.000 1.680 ;
        RECT  2.780 1.440 4.000 1.680 ;
        RECT  7.170 1.130 7.410 1.970 ;
        RECT  2.230 3.260 2.470 3.810 ;
        RECT  7.390 1.730 7.630 3.810 ;
        RECT  2.230 3.570 7.630 3.810 ;
        RECT  8.640 1.440 8.890 3.230 ;
        RECT  9.820 2.190 10.060 2.870 ;
        RECT  9.560 2.630 10.060 2.870 ;
        RECT  7.900 1.440 8.150 3.720 ;
        RECT  9.560 2.630 9.800 3.720 ;
        RECT  7.900 3.480 9.800 3.720 ;
        RECT  10.030 1.440 10.540 1.920 ;
        RECT  9.130 1.680 10.540 1.920 ;
        RECT  9.130 1.680 9.370 2.480 ;
        RECT  10.300 1.440 10.540 3.510 ;
        RECT  10.040 3.110 10.540 3.510 ;
        RECT  11.370 1.520 11.940 1.760 ;
        RECT  11.370 1.520 11.610 3.370 ;
        RECT  11.370 3.130 11.920 3.370 ;
        RECT  12.910 1.640 13.310 2.040 ;
        RECT  12.370 1.720 13.310 2.040 ;
        RECT  12.370 1.720 12.610 2.300 ;
        RECT  11.880 2.060 12.610 2.300 ;
        RECT  11.880 2.060 12.120 2.640 ;
        RECT  13.560 2.350 13.800 2.900 ;
        RECT  13.070 2.660 13.800 2.900 ;
        RECT  13.070 1.640 13.310 3.580 ;
        RECT  12.930 3.360 13.170 3.890 ;
        RECT  14.830 2.490 15.650 2.730 ;
        RECT  12.560 2.600 12.800 3.150 ;
        RECT  10.860 1.440 11.110 3.930 ;
        RECT  10.860 3.690 12.690 3.930 ;
        RECT  12.450 2.910 12.690 4.370 ;
        RECT  14.830 2.490 15.070 4.370 ;
        RECT  12.450 4.130 15.070 4.370 ;
    END
END sdnfb2

MACRO sdnfb1
    CLASS CORE ;
    FOREIGN sdnfb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.451  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.210 2.230 5.610 2.720 ;
        RECT  5.100 2.020 5.540 2.460 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.020 4.520 2.460 ;
        RECT  4.120 1.890 4.520 2.460 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.384  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.580 1.460 14.500 1.900 ;
        RECT  13.580 1.150 14.020 1.900 ;
        RECT  13.580 1.150 13.980 3.410 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.228  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.180 2.580 15.550 3.020 ;
        RECT  15.310 1.110 15.550 3.020 ;
        RECT  15.210 2.580 15.450 3.900 ;
        RECT  15.130 1.110 15.550 1.530 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.390 2.520 0.790 2.920 ;
        RECT  0.130 2.580 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.290 2.450 2.740 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.680 5.600 ;
        RECT  14.480 4.610 14.880 5.600 ;
        RECT  12.180 4.610 12.580 5.600 ;
        RECT  9.380 3.960 9.620 5.600 ;
        RECT  5.730 4.180 5.970 5.600 ;
        RECT  3.180 4.360 3.580 5.600 ;
        RECT  0.800 4.570 1.200 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.680 0.740 ;
        RECT  14.390 0.000 14.790 1.220 ;
        RECT  12.240 0.000 12.640 0.890 ;
        RECT  9.390 0.000 9.630 1.440 ;
        RECT  6.610 0.000 7.010 0.890 ;
        RECT  3.260 0.000 3.500 1.200 ;
        RECT  0.820 0.000 1.060 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.270 2.090 ;
        RECT  1.030 1.850 1.270 3.530 ;
        RECT  1.030 2.560 1.480 2.960 ;
        RECT  1.030 2.560 1.280 3.530 ;
        RECT  0.150 3.290 1.280 3.530 ;
        RECT  1.510 1.770 1.910 2.170 ;
        RECT  1.510 1.930 3.590 2.170 ;
        RECT  3.190 1.930 3.590 2.370 ;
        RECT  1.720 1.930 1.960 3.440 ;
        RECT  1.530 3.200 1.770 3.750 ;
        RECT  5.020 1.540 6.090 1.780 ;
        RECT  5.850 2.230 6.410 2.630 ;
        RECT  5.850 1.540 6.090 3.320 ;
        RECT  5.080 3.080 6.090 3.320 ;
        RECT  6.380 1.640 6.930 1.890 ;
        RECT  6.690 1.640 6.930 2.360 ;
        RECT  6.770 2.110 7.010 3.230 ;
        RECT  6.380 2.990 7.010 3.230 ;
        RECT  1.980 0.980 3.020 1.220 ;
        RECT  3.760 0.980 4.930 1.220 ;
        RECT  4.690 1.060 6.440 1.300 ;
        RECT  6.270 1.130 7.410 1.370 ;
        RECT  2.780 0.980 3.020 1.680 ;
        RECT  3.760 0.980 4.000 1.680 ;
        RECT  2.780 1.440 4.000 1.680 ;
        RECT  7.170 1.130 7.410 1.840 ;
        RECT  2.230 3.260 2.470 3.810 ;
        RECT  7.400 1.600 7.640 3.810 ;
        RECT  2.230 3.570 7.640 3.810 ;
        RECT  8.640 1.290 8.890 3.230 ;
        RECT  9.810 2.190 10.050 2.860 ;
        RECT  9.560 2.620 10.050 2.860 ;
        RECT  7.900 1.290 8.150 3.720 ;
        RECT  9.560 2.620 9.800 3.720 ;
        RECT  7.900 3.480 9.800 3.720 ;
        RECT  10.040 1.440 10.450 1.920 ;
        RECT  9.130 1.680 10.530 1.920 ;
        RECT  9.130 1.680 9.370 2.470 ;
        RECT  10.290 1.680 10.530 3.510 ;
        RECT  10.040 3.110 10.530 3.510 ;
        RECT  11.370 1.520 11.940 1.760 ;
        RECT  11.370 1.520 11.610 3.370 ;
        RECT  11.370 3.130 11.920 3.370 ;
        RECT  12.370 1.720 13.310 1.960 ;
        RECT  12.910 1.640 13.310 2.040 ;
        RECT  12.370 1.720 12.610 2.300 ;
        RECT  11.880 2.060 12.610 2.300 ;
        RECT  11.880 2.060 12.120 2.640 ;
        RECT  13.070 1.640 13.310 3.890 ;
        RECT  12.850 3.400 13.310 3.890 ;
        RECT  14.220 2.520 14.460 3.890 ;
        RECT  12.850 3.650 14.460 3.890 ;
        RECT  14.820 1.830 15.060 2.370 ;
        RECT  12.560 2.600 12.800 3.150 ;
        RECT  10.860 1.440 11.110 3.930 ;
        RECT  10.860 3.690 12.610 3.930 ;
        RECT  12.370 2.910 12.610 4.370 ;
        RECT  14.700 2.140 14.940 4.370 ;
        RECT  12.370 4.130 14.940 4.370 ;
    END
END sdnfb1

MACRO sdcrq4
    CLASS CORE ;
    FOREIGN sdcrq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.392  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.580 2.500 10.020 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.320 2.340 5.730 2.740 ;
        RECT  5.100 2.020 5.540 2.460 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.300 2.820 ;
        RECT  4.060 2.050 4.300 2.820 ;
        RECT  3.420 2.580 3.860 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.844  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.320 3.940 17.800 4.340 ;
        RECT  17.370 1.530 17.800 4.340 ;
        RECT  15.380 1.530 17.800 1.930 ;
        RECT  14.650 1.310 15.620 1.550 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.520 0.800 2.920 ;
        RECT  0.130 2.520 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.290 2.450 2.740 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.920 5.600 ;
        RECT  17.370 4.620 17.770 5.600 ;
        RECT  16.060 4.620 16.460 5.600 ;
        RECT  14.750 4.620 15.150 5.600 ;
        RECT  13.340 4.300 13.580 5.600 ;
        RECT  10.420 4.710 10.820 5.600 ;
        RECT  9.150 4.710 9.550 5.600 ;
        RECT  5.810 4.180 6.050 5.600 ;
        RECT  3.260 4.360 3.500 5.600 ;
        RECT  0.880 4.510 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.920 0.740 ;
        RECT  16.690 0.000 17.090 0.890 ;
        RECT  15.330 0.000 15.730 0.890 ;
        RECT  12.800 0.000 13.040 1.420 ;
        RECT  9.840 0.000 10.080 1.640 ;
        RECT  7.320 0.000 7.720 0.890 ;
        RECT  3.260 0.000 3.500 1.200 ;
        RECT  0.820 0.000 1.060 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.280 2.090 ;
        RECT  1.040 2.560 1.480 2.960 ;
        RECT  1.040 1.850 1.280 3.530 ;
        RECT  0.150 3.290 1.280 3.530 ;
        RECT  1.590 1.660 1.830 2.210 ;
        RECT  1.590 1.970 3.510 2.210 ;
        RECT  1.720 1.970 1.960 3.440 ;
        RECT  1.530 3.200 1.770 3.750 ;
        RECT  5.020 1.540 6.020 1.780 ;
        RECT  5.780 1.540 6.020 2.100 ;
        RECT  5.970 2.340 6.410 2.740 ;
        RECT  5.970 1.860 6.210 3.320 ;
        RECT  5.080 3.080 6.210 3.320 ;
        RECT  1.980 0.980 3.020 1.220 ;
        RECT  4.230 0.980 7.090 1.220 ;
        RECT  6.860 1.130 7.400 1.370 ;
        RECT  2.780 0.980 3.020 1.700 ;
        RECT  4.230 0.980 4.470 1.700 ;
        RECT  2.780 1.460 4.780 1.700 ;
        RECT  7.160 1.130 7.400 1.880 ;
        RECT  2.230 3.260 2.470 3.840 ;
        RECT  7.390 1.640 7.630 3.700 ;
        RECT  7.080 3.460 7.630 3.700 ;
        RECT  2.230 3.600 4.780 3.840 ;
        RECT  4.540 1.460 4.780 4.000 ;
        RECT  4.380 3.600 4.780 4.000 ;
        RECT  8.380 1.460 8.960 1.700 ;
        RECT  8.380 1.460 8.620 3.990 ;
        RECT  8.380 3.750 10.320 3.990 ;
        RECT  7.960 0.980 9.600 1.220 ;
        RECT  9.360 0.980 9.600 2.120 ;
        RECT  9.360 1.880 10.500 2.120 ;
        RECT  10.260 1.880 10.500 2.820 ;
        RECT  10.260 2.410 10.700 2.820 ;
        RECT  7.900 1.050 8.140 3.390 ;
        RECT  10.500 1.240 10.990 1.640 ;
        RECT  10.750 1.240 10.990 2.020 ;
        RECT  10.750 1.780 11.250 2.020 ;
        RECT  8.890 2.270 9.130 3.510 ;
        RECT  11.010 1.780 11.250 3.510 ;
        RECT  8.890 3.270 11.590 3.510 ;
        RECT  6.460 1.550 6.700 2.100 ;
        RECT  6.650 1.860 6.890 2.630 ;
        RECT  6.650 2.230 7.100 2.630 ;
        RECT  6.770 2.230 7.010 3.230 ;
        RECT  6.460 2.990 7.010 3.230 ;
        RECT  6.460 2.990 6.700 4.470 ;
        RECT  6.460 4.230 12.540 4.470 ;
        RECT  12.060 1.220 12.300 2.420 ;
        RECT  12.060 2.180 12.730 2.420 ;
        RECT  12.490 2.180 12.730 3.430 ;
        RECT  12.490 3.190 13.070 3.430 ;
        RECT  11.240 1.300 11.800 1.540 ;
        RECT  11.560 1.300 11.800 2.900 ;
        RECT  11.560 2.660 12.250 2.900 ;
        RECT  14.190 2.280 14.430 3.100 ;
        RECT  13.480 2.860 14.430 3.100 ;
        RECT  13.480 2.860 13.720 3.430 ;
        RECT  12.010 2.660 12.250 3.910 ;
        RECT  13.310 3.190 13.550 3.910 ;
        RECT  12.010 3.670 13.550 3.910 ;
        RECT  13.420 1.070 14.320 1.310 ;
        RECT  13.420 1.070 13.660 2.040 ;
        RECT  13.000 1.800 14.910 2.040 ;
        RECT  14.670 2.390 17.120 2.790 ;
        RECT  13.000 1.800 13.240 2.930 ;
        RECT  14.670 1.800 14.910 3.800 ;
        RECT  13.970 3.560 14.910 3.800 ;
    END
END sdcrq4

MACRO sdcrq2
    CLASS CORE ;
    FOREIGN sdcrq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.412  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.300 2.580 16.740 3.020 ;
        RECT  15.950 2.350 16.350 2.820 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.504  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.790 3.400 17.800 3.640 ;
        RECT  17.490 1.210 17.800 3.640 ;
        RECT  17.420 1.210 17.800 1.900 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.920 5.600 ;
        RECT  17.450 4.170 17.690 5.600 ;
        RECT  16.150 3.950 16.390 5.600 ;
        RECT  14.830 3.960 15.070 5.600 ;
        RECT  11.810 4.350 12.050 5.600 ;
        RECT  10.450 4.350 10.690 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.920 0.740 ;
        RECT  16.060 0.000 16.480 0.890 ;
        RECT  14.310 0.000 14.710 0.890 ;
        RECT  11.530 0.000 11.770 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.550 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.060 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.060 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.510 4.110 ;
        RECT  10.320 1.750 10.560 3.630 ;
        RECT  10.320 3.130 10.660 3.630 ;
        RECT  10.320 3.390 11.540 3.630 ;
        RECT  9.580 1.270 11.060 1.510 ;
        RECT  10.820 1.270 11.060 2.600 ;
        RECT  10.820 2.360 12.320 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  12.230 1.830 12.810 2.070 ;
        RECT  12.570 1.830 12.810 3.100 ;
        RECT  11.300 2.860 12.810 3.100 ;
        RECT  12.330 2.860 12.570 3.630 ;
        RECT  12.330 3.390 12.900 3.630 ;
        RECT  9.850 3.870 12.530 4.110 ;
        RECT  12.290 3.870 12.530 4.620 ;
        RECT  12.290 4.380 13.260 4.620 ;
        RECT  13.800 1.610 14.050 2.010 ;
        RECT  13.800 1.610 14.040 3.960 ;
        RECT  13.800 3.720 14.380 3.960 ;
        RECT  13.050 1.130 15.230 1.370 ;
        RECT  13.050 1.130 13.290 3.180 ;
        RECT  14.990 1.130 15.230 2.960 ;
        RECT  13.050 2.940 13.560 3.180 ;
        RECT  13.320 2.940 13.560 3.710 ;
        RECT  15.620 1.420 15.860 2.110 ;
        RECT  15.470 1.870 16.840 2.110 ;
        RECT  16.600 2.100 17.220 2.340 ;
        RECT  16.980 2.100 17.220 2.710 ;
        RECT  14.280 2.770 14.520 3.480 ;
        RECT  15.470 1.870 15.710 3.710 ;
        RECT  14.280 3.240 15.710 3.480 ;
        RECT  15.330 3.300 15.730 3.710 ;
    END
END sdcrq2

MACRO sdcrq1
    CLASS CORE ;
    FOREIGN sdcrq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.412  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.300 2.580 16.740 3.020 ;
        RECT  15.950 2.350 16.350 2.820 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.252  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.860 3.400 17.240 4.140 ;
        RECT  16.980 1.140 17.240 4.140 ;
        RECT  16.780 1.140 17.240 1.460 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.360 5.600 ;
        RECT  16.150 3.950 16.390 5.600 ;
        RECT  14.830 3.960 15.070 5.600 ;
        RECT  11.810 4.350 12.050 5.600 ;
        RECT  10.450 4.350 10.690 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.360 0.740 ;
        RECT  16.030 0.000 16.450 0.980 ;
        RECT  14.280 0.000 14.680 0.890 ;
        RECT  11.530 0.000 11.770 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.550 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.150 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.150 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.510 4.110 ;
        RECT  10.320 1.750 10.560 3.630 ;
        RECT  10.320 3.130 10.660 3.630 ;
        RECT  10.320 3.390 11.540 3.630 ;
        RECT  9.580 1.270 11.060 1.510 ;
        RECT  10.820 1.270 11.060 2.600 ;
        RECT  10.820 2.360 12.320 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  12.230 1.830 12.810 2.070 ;
        RECT  12.570 1.830 12.810 3.100 ;
        RECT  11.300 2.860 12.810 3.100 ;
        RECT  12.330 2.860 12.570 3.630 ;
        RECT  12.330 3.390 12.900 3.630 ;
        RECT  9.850 3.870 12.530 4.110 ;
        RECT  12.290 3.870 12.530 4.620 ;
        RECT  12.290 4.380 13.260 4.620 ;
        RECT  13.790 1.610 14.040 2.010 ;
        RECT  13.800 1.610 14.040 3.960 ;
        RECT  13.800 3.720 14.380 3.960 ;
        RECT  13.050 1.130 15.230 1.370 ;
        RECT  13.050 1.130 13.290 3.180 ;
        RECT  14.990 1.130 15.230 2.960 ;
        RECT  13.050 2.940 13.560 3.180 ;
        RECT  13.320 2.940 13.560 3.710 ;
        RECT  15.590 1.420 15.830 1.990 ;
        RECT  15.470 1.750 16.690 1.990 ;
        RECT  14.280 2.770 14.520 3.480 ;
        RECT  15.470 1.750 15.710 3.710 ;
        RECT  14.280 3.240 15.710 3.480 ;
        RECT  15.330 3.300 15.730 3.710 ;
    END
END sdcrq1

MACRO sdcrn4
    CLASS CORE ;
    FOREIGN sdcrn4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.580 7.510 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.040 1.680 14.500 2.460 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.453  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.600 2.820 3.020 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.876  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.410 1.530 17.130 1.930 ;
        RECT  16.890 1.110 17.130 1.930 ;
        RECT  16.270 1.530 16.710 3.020 ;
        RECT  16.250 3.820 16.650 4.140 ;
        RECT  16.270 1.530 16.650 4.140 ;
        RECT  14.910 3.820 16.650 4.060 ;
        RECT  15.410 1.110 15.650 1.930 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.670 3.070 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.210 3.020 ;
        RECT  3.970 2.210 4.210 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.360 5.600 ;
        RECT  15.680 4.420 16.080 5.600 ;
        RECT  14.340 4.420 14.740 5.600 ;
        RECT  12.300 4.710 12.700 5.600 ;
        RECT  10.900 4.710 11.300 5.600 ;
        RECT  8.060 4.710 8.460 5.600 ;
        RECT  6.740 4.710 7.130 5.600 ;
        RECT  3.260 4.520 3.660 5.600 ;
        RECT  0.780 4.620 1.180 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.360 0.740 ;
        RECT  16.070 0.000 16.470 0.980 ;
        RECT  14.590 0.000 14.990 0.980 ;
        RECT  12.980 0.000 13.380 0.890 ;
        RECT  7.290 0.000 7.530 1.650 ;
        RECT  3.180 1.080 3.800 1.320 ;
        RECT  3.560 0.000 3.800 1.320 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.340 1.820 ;
        RECT  1.100 1.580 1.340 2.910 ;
        RECT  1.000 2.700 1.240 3.590 ;
        RECT  0.150 3.350 1.240 3.590 ;
        RECT  1.590 2.100 3.510 2.340 ;
        RECT  1.590 1.760 1.830 3.230 ;
        RECT  1.530 3.070 1.770 3.670 ;
        RECT  1.980 0.980 2.770 1.220 ;
        RECT  2.530 0.980 2.770 1.860 ;
        RECT  2.530 1.620 4.700 1.860 ;
        RECT  4.460 1.070 4.700 3.650 ;
        RECT  2.150 3.330 4.790 3.570 ;
        RECT  4.460 3.250 4.790 3.650 ;
        RECT  4.450 3.330 4.790 3.650 ;
        RECT  5.710 1.540 6.290 1.780 ;
        RECT  5.710 1.540 5.950 2.270 ;
        RECT  5.700 2.190 5.940 3.510 ;
        RECT  5.700 3.270 7.790 3.510 ;
        RECT  5.220 1.420 5.470 1.740 ;
        RECT  5.220 1.420 5.460 4.140 ;
        RECT  5.140 3.740 5.460 4.140 ;
        RECT  8.030 2.640 8.270 3.990 ;
        RECT  5.140 3.750 8.270 3.990 ;
        RECT  5.140 3.750 5.540 4.140 ;
        RECT  6.240 2.060 8.300 2.300 ;
        RECT  8.060 1.440 8.300 2.300 ;
        RECT  8.090 2.160 8.750 2.400 ;
        RECT  6.240 2.060 6.480 2.650 ;
        RECT  8.510 2.160 8.750 3.090 ;
        RECT  8.740 2.850 8.980 3.610 ;
        RECT  9.480 1.510 10.230 1.750 ;
        RECT  9.990 1.510 10.230 3.510 ;
        RECT  9.990 3.260 10.570 3.510 ;
        RECT  8.740 1.480 9.230 1.880 ;
        RECT  8.990 1.480 9.230 2.610 ;
        RECT  8.990 2.370 9.750 2.610 ;
        RECT  11.630 2.190 11.870 2.800 ;
        RECT  11.070 2.560 11.870 2.800 ;
        RECT  11.070 2.560 11.310 3.450 ;
        RECT  9.510 2.370 9.750 3.990 ;
        RECT  11.000 3.220 11.240 3.990 ;
        RECT  9.510 3.750 11.240 3.990 ;
        RECT  10.500 1.520 12.320 1.760 ;
        RECT  10.500 1.520 10.740 3.020 ;
        RECT  12.120 1.610 12.360 3.990 ;
        RECT  11.480 3.730 12.360 3.990 ;
        RECT  8.500 0.980 12.740 1.220 ;
        RECT  12.510 1.130 13.320 1.370 ;
        RECT  13.080 1.130 13.320 3.580 ;
        RECT  13.560 1.070 14.210 1.310 ;
        RECT  13.560 1.070 13.800 3.780 ;
        RECT  12.600 2.620 12.840 4.470 ;
        RECT  5.970 4.230 13.920 4.470 ;
        RECT  13.680 3.500 13.920 4.470 ;
        RECT  5.490 4.380 6.240 4.620 ;
    END
END sdcrn4

MACRO sdcrn2
    CLASS CORE ;
    FOREIGN sdcrn2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.412  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.300 2.580 16.740 3.020 ;
        RECT  15.950 2.310 16.350 2.820 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.504  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.860 1.460 17.300 1.900 ;
        RECT  16.790 3.400 17.220 3.720 ;
        RECT  16.980 1.460 17.220 3.720 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.920 5.600 ;
        RECT  17.450 4.170 17.690 5.600 ;
        RECT  16.150 3.950 16.390 5.600 ;
        RECT  14.830 3.960 15.070 5.600 ;
        RECT  11.810 4.350 12.050 5.600 ;
        RECT  10.450 4.350 10.690 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.920 0.740 ;
        RECT  16.060 0.000 16.480 0.890 ;
        RECT  14.310 0.000 14.710 0.890 ;
        RECT  11.530 0.000 11.770 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.560 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.150 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.150 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.510 4.110 ;
        RECT  10.320 1.750 10.560 3.630 ;
        RECT  10.320 3.130 10.660 3.630 ;
        RECT  10.320 3.390 11.540 3.630 ;
        RECT  9.580 1.270 11.060 1.510 ;
        RECT  10.820 1.270 11.060 2.600 ;
        RECT  10.820 2.360 12.320 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  12.230 1.830 12.810 2.070 ;
        RECT  12.570 1.830 12.810 3.100 ;
        RECT  11.300 2.860 12.810 3.100 ;
        RECT  12.330 2.860 12.570 3.630 ;
        RECT  12.330 3.390 12.900 3.630 ;
        RECT  9.850 3.870 12.530 4.110 ;
        RECT  12.290 3.870 12.530 4.620 ;
        RECT  12.290 4.380 13.260 4.620 ;
        RECT  13.800 1.610 14.050 2.010 ;
        RECT  13.800 1.610 14.040 3.960 ;
        RECT  13.800 3.720 14.380 3.960 ;
        RECT  13.050 1.130 15.230 1.370 ;
        RECT  13.050 1.130 13.290 3.180 ;
        RECT  14.990 1.130 15.230 2.960 ;
        RECT  13.050 2.940 13.560 3.180 ;
        RECT  13.320 2.940 13.560 3.710 ;
        RECT  15.620 1.420 15.860 1.980 ;
        RECT  14.280 2.770 14.520 3.480 ;
        RECT  15.470 1.740 15.710 3.710 ;
        RECT  14.280 3.240 15.710 3.480 ;
        RECT  15.330 3.300 15.730 3.710 ;
    END
END sdcrn2

MACRO sdcrn1
    CLASS CORE ;
    FOREIGN sdcrn1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.412  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.300 2.580 16.740 3.020 ;
        RECT  15.950 2.310 16.350 2.820 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.276  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.790 3.400 17.230 3.720 ;
        RECT  16.980 1.460 17.230 3.720 ;
        RECT  16.830 1.190 17.100 1.900 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.360 5.600 ;
        RECT  16.150 3.950 16.390 5.600 ;
        RECT  14.830 3.960 15.070 5.600 ;
        RECT  11.810 4.350 12.050 5.600 ;
        RECT  10.450 4.350 10.690 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.360 0.740 ;
        RECT  16.030 0.000 16.450 0.980 ;
        RECT  14.280 0.000 14.680 0.890 ;
        RECT  11.530 0.000 11.770 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.550 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.150 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.150 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.510 4.110 ;
        RECT  10.320 1.750 10.560 3.630 ;
        RECT  10.320 3.130 10.660 3.630 ;
        RECT  10.320 3.390 11.540 3.630 ;
        RECT  9.580 1.270 11.060 1.510 ;
        RECT  10.820 1.270 11.060 2.600 ;
        RECT  10.820 2.360 12.320 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  12.230 1.830 12.810 2.070 ;
        RECT  12.570 1.830 12.810 3.100 ;
        RECT  11.300 2.860 12.810 3.100 ;
        RECT  12.330 2.860 12.570 3.630 ;
        RECT  12.330 3.390 12.900 3.630 ;
        RECT  9.850 3.870 12.530 4.110 ;
        RECT  12.290 3.870 12.530 4.620 ;
        RECT  12.290 4.380 13.260 4.620 ;
        RECT  13.790 1.610 14.040 2.010 ;
        RECT  13.800 1.610 14.040 3.960 ;
        RECT  13.800 3.720 14.380 3.960 ;
        RECT  13.050 1.130 15.230 1.370 ;
        RECT  13.050 1.130 13.290 3.180 ;
        RECT  14.990 1.130 15.230 2.960 ;
        RECT  13.050 2.940 13.560 3.180 ;
        RECT  13.320 2.940 13.560 3.710 ;
        RECT  15.590 1.420 15.830 1.980 ;
        RECT  14.280 2.770 14.520 3.480 ;
        RECT  15.470 1.740 15.710 3.710 ;
        RECT  14.280 3.240 15.710 3.480 ;
        RECT  15.330 3.300 15.730 3.710 ;
    END
END sdcrn1

MACRO sdcrb4
    CLASS CORE ;
    FOREIGN sdcrb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.690 1.750 17.300 2.540 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.580 5.540 3.020 ;
        RECT  4.980 2.770 5.380 3.170 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.340 2.480 3.860 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.944  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.380 1.220 15.270 1.460 ;
        RECT  13.710 3.190 15.260 3.430 ;
        RECT  15.020 2.800 15.260 3.430 ;
        RECT  13.710 1.220 13.950 3.430 ;
        RECT  12.940 2.020 13.950 2.460 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.080  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.650 2.020 19.510 2.460 ;
        RECT  19.110 1.060 19.510 2.460 ;
        RECT  18.790 2.020 19.190 4.240 ;
        RECT  17.650 2.020 18.050 2.900 ;
        RECT  17.620 1.050 18.020 2.280 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.800 2.830 ;
        RECT  0.120 2.430 0.500 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.870 4.220 2.110 ;
        RECT  2.470 1.870 2.870 2.570 ;
        RECT  2.300 2.570 2.740 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.160 5.600 ;
        RECT  19.610 4.480 20.010 5.600 ;
        RECT  18.300 3.170 18.540 5.600 ;
        RECT  16.900 4.360 17.300 5.600 ;
        RECT  15.510 4.360 15.910 5.600 ;
        RECT  14.200 4.360 14.600 5.600 ;
        RECT  12.890 4.360 13.290 5.600 ;
        RECT  10.110 4.400 10.510 5.600 ;
        RECT  8.840 4.110 9.240 5.600 ;
        RECT  5.490 4.550 5.890 5.600 ;
        RECT  4.220 4.620 4.620 5.600 ;
        RECT  1.990 4.620 2.390 5.600 ;
        RECT  0.720 4.550 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.160 0.740 ;
        RECT  18.370 0.000 18.770 0.980 ;
        RECT  16.770 0.000 17.170 1.220 ;
        RECT  14.130 0.000 14.530 0.980 ;
        RECT  12.650 0.000 13.050 0.980 ;
        RECT  9.360 0.000 9.760 1.770 ;
        RECT  5.230 0.000 5.630 1.060 ;
        RECT  4.530 0.000 4.930 0.990 ;
        RECT  0.740 0.000 1.140 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.500 0.470 2.190 ;
        RECT  0.230 1.950 1.280 2.190 ;
        RECT  1.040 2.420 1.480 2.820 ;
        RECT  1.040 1.950 1.280 3.580 ;
        RECT  0.150 3.340 1.280 3.580 ;
        RECT  1.590 1.490 1.830 2.200 ;
        RECT  4.120 2.650 4.520 3.050 ;
        RECT  4.120 2.650 4.360 3.500 ;
        RECT  1.720 3.260 4.360 3.500 ;
        RECT  1.720 1.960 1.960 4.340 ;
        RECT  1.460 3.940 1.960 4.340 ;
        RECT  4.780 1.790 5.410 2.030 ;
        RECT  5.170 1.790 5.410 2.310 ;
        RECT  5.170 2.070 6.080 2.310 ;
        RECT  5.840 2.070 6.080 3.060 ;
        RECT  5.780 2.820 6.020 3.730 ;
        RECT  4.920 3.490 6.020 3.730 ;
        RECT  6.400 2.470 6.840 2.870 ;
        RECT  6.400 1.760 6.640 3.380 ;
        RECT  6.310 3.140 6.550 3.700 ;
        RECT  5.880 1.060 7.230 1.300 ;
        RECT  3.240 1.090 3.640 1.550 ;
        RECT  5.880 1.060 6.120 1.550 ;
        RECT  3.240 1.310 6.120 1.550 ;
        RECT  6.990 1.060 7.230 1.960 ;
        RECT  3.190 3.740 4.670 3.980 ;
        RECT  4.430 3.970 6.600 4.210 ;
        RECT  6.360 3.970 6.600 4.620 ;
        RECT  7.080 1.720 7.320 4.620 ;
        RECT  6.360 4.380 7.320 4.620 ;
        RECT  8.200 1.810 8.450 2.410 ;
        RECT  8.040 2.170 8.280 3.890 ;
        RECT  8.040 3.490 9.810 3.730 ;
        RECT  8.040 3.490 8.470 3.890 ;
        RECT  7.470 0.980 7.710 1.530 ;
        RECT  7.470 1.290 9.040 1.530 ;
        RECT  8.800 1.290 9.040 2.250 ;
        RECT  8.800 2.010 9.620 2.250 ;
        RECT  9.380 2.010 9.620 2.550 ;
        RECT  9.380 2.310 9.960 2.550 ;
        RECT  7.560 1.290 7.800 4.280 ;
        RECT  7.580 4.040 7.820 4.620 ;
        RECT  10.180 1.420 10.420 2.030 ;
        RECT  8.520 2.670 8.760 3.250 ;
        RECT  8.520 3.010 10.440 3.250 ;
        RECT  10.200 1.790 10.440 3.960 ;
        RECT  10.200 3.720 11.080 3.960 ;
        RECT  11.410 1.480 11.650 3.000 ;
        RECT  11.650 0.990 12.350 1.230 ;
        RECT  12.110 0.990 12.350 3.520 ;
        RECT  12.110 3.280 12.740 3.520 ;
        RECT  15.650 1.050 15.890 2.030 ;
        RECT  14.200 1.880 15.850 2.280 ;
        RECT  15.610 1.790 15.850 3.640 ;
        RECT  15.600 3.400 16.680 3.640 ;
        RECT  10.680 0.990 11.270 1.230 ;
        RECT  16.090 2.270 16.330 3.150 ;
        RECT  16.090 2.910 17.250 3.150 ;
        RECT  10.680 0.990 10.920 3.480 ;
        RECT  10.680 3.240 11.770 3.480 ;
        RECT  11.530 3.240 11.770 4.120 ;
        RECT  17.010 2.910 17.250 4.120 ;
        RECT  11.530 3.880 17.250 4.120 ;
    END
END sdcrb4

MACRO sdcrb2
    CLASS CORE ;
    FOREIGN sdcrb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.700 2.580 16.180 3.020 ;
        RECT  15.700 2.310 15.940 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.222  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.300 3.050 18.980 3.580 ;
        RECT  18.740 1.650 18.980 3.580 ;
        RECT  18.380 1.650 18.980 1.890 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.232  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.860 1.460 17.300 1.900 ;
        RECT  17.000 1.460 17.240 2.870 ;
        RECT  16.920 2.660 17.160 3.450 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.290 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.600 5.600 ;
        RECT  19.010 4.170 19.250 5.600 ;
        RECT  17.590 4.170 17.830 5.600 ;
        RECT  16.240 4.170 16.480 5.600 ;
        RECT  14.830 4.160 15.070 5.600 ;
        RECT  11.810 4.350 12.050 5.600 ;
        RECT  10.450 4.350 10.690 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.600 0.740 ;
        RECT  19.130 0.000 19.370 1.400 ;
        RECT  17.710 0.000 17.950 1.400 ;
        RECT  16.330 0.000 16.570 1.400 ;
        RECT  14.310 0.000 14.710 0.890 ;
        RECT  11.530 0.000 11.770 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.550 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.150 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.150 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.510 4.110 ;
        RECT  10.320 1.750 10.560 3.630 ;
        RECT  10.320 3.130 10.660 3.630 ;
        RECT  10.320 3.390 11.540 3.630 ;
        RECT  9.580 1.270 11.060 1.510 ;
        RECT  10.820 1.270 11.060 2.600 ;
        RECT  10.820 2.360 12.320 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  12.230 1.830 12.810 2.070 ;
        RECT  12.570 1.830 12.810 3.100 ;
        RECT  11.300 2.860 12.810 3.100 ;
        RECT  12.330 2.860 12.570 3.630 ;
        RECT  12.330 3.390 12.900 3.630 ;
        RECT  9.850 3.870 12.530 4.110 ;
        RECT  12.290 3.870 12.530 4.490 ;
        RECT  12.290 4.250 13.260 4.490 ;
        RECT  13.800 1.610 14.050 2.010 ;
        RECT  13.800 1.610 14.040 3.960 ;
        RECT  13.800 3.720 14.380 3.960 ;
        RECT  13.050 1.130 15.000 1.370 ;
        RECT  14.760 1.130 15.000 2.800 ;
        RECT  13.050 1.130 13.290 3.180 ;
        RECT  14.910 2.560 15.310 2.960 ;
        RECT  13.050 2.940 13.560 3.180 ;
        RECT  13.320 2.940 13.560 3.710 ;
        RECT  15.620 1.420 15.860 1.980 ;
        RECT  15.620 1.740 16.600 1.980 ;
        RECT  16.360 1.740 16.600 2.350 ;
        RECT  17.520 2.180 18.450 2.420 ;
        RECT  14.280 2.770 14.520 3.480 ;
        RECT  14.280 3.240 15.240 3.480 ;
        RECT  15.000 3.260 15.730 3.500 ;
        RECT  15.330 3.260 15.730 3.750 ;
        RECT  16.420 2.110 16.660 3.930 ;
        RECT  15.330 3.510 16.660 3.750 ;
        RECT  17.520 2.180 17.760 3.930 ;
        RECT  16.420 3.690 17.760 3.930 ;
    END
END sdcrb2

MACRO sdcrb1
    CLASS CORE ;
    FOREIGN sdcrb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.300 3.700 16.740 4.140 ;
        RECT  16.030 3.700 16.740 3.940 ;
        RECT  16.030 2.880 16.270 3.940 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.060  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.620 1.460 17.300 1.900 ;
        RECT  16.620 3.130 17.180 3.370 ;
        RECT  16.940 1.460 17.180 3.370 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.049  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.980 2.580 18.360 3.020 ;
        RECT  17.980 1.570 18.250 3.450 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 18.480 5.600 ;
        RECT  17.270 4.020 17.510 5.600 ;
        RECT  16.100 4.710 16.500 5.600 ;
        RECT  14.830 4.160 15.070 5.600 ;
        RECT  11.810 4.350 12.050 5.600 ;
        RECT  10.450 4.350 10.690 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 18.480 0.740 ;
        RECT  17.420 0.000 17.660 1.230 ;
        RECT  14.310 0.000 14.710 0.890 ;
        RECT  11.530 0.000 11.770 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.550 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.150 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.150 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.510 4.110 ;
        RECT  10.320 1.750 10.560 3.630 ;
        RECT  10.320 3.130 10.740 3.630 ;
        RECT  10.320 3.390 11.540 3.630 ;
        RECT  9.580 1.270 11.060 1.510 ;
        RECT  10.820 1.270 11.060 2.600 ;
        RECT  10.820 2.360 12.320 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  12.230 1.830 12.810 2.070 ;
        RECT  12.570 1.830 12.810 3.100 ;
        RECT  11.300 2.860 12.810 3.100 ;
        RECT  12.330 2.860 12.570 3.630 ;
        RECT  12.330 3.390 12.900 3.630 ;
        RECT  9.850 3.870 12.530 4.110 ;
        RECT  12.290 3.870 12.530 4.490 ;
        RECT  12.290 4.250 13.260 4.490 ;
        RECT  13.800 1.610 14.050 2.010 ;
        RECT  13.800 1.610 14.040 3.960 ;
        RECT  13.800 3.720 14.380 3.960 ;
        RECT  13.050 1.130 15.230 1.370 ;
        RECT  13.050 1.130 13.290 3.180 ;
        RECT  14.990 1.130 15.230 2.960 ;
        RECT  13.050 2.940 13.560 3.180 ;
        RECT  13.320 2.940 13.560 3.710 ;
        RECT  15.620 1.420 15.860 2.420 ;
        RECT  15.490 2.180 16.680 2.420 ;
        RECT  16.280 2.180 16.680 2.580 ;
        RECT  14.280 2.770 14.520 3.480 ;
        RECT  15.490 2.180 15.730 3.480 ;
        RECT  14.280 3.240 15.730 3.480 ;
        RECT  15.410 3.240 15.650 3.810 ;
    END
END sdcrb1

MACRO sdcfq4
    CLASS CORE ;
    FOREIGN sdcfq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.818  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.770 3.020 14.170 3.420 ;
        RECT  13.500 3.370 14.050 3.610 ;
        RECT  13.500 3.370 13.740 4.380 ;
        RECT  12.670 4.140 13.740 4.380 ;
        RECT  11.300 4.380 12.910 4.620 ;
        RECT  11.300 3.350 11.540 4.620 ;
        RECT  10.390 3.350 11.540 3.590 ;
        RECT  10.390 2.870 10.630 3.590 ;
        RECT  9.580 2.870 10.630 3.120 ;
        RECT  9.580 2.560 10.070 3.120 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.441  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.010 2.130 5.540 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.540 2.020 4.420 2.460 ;
        RECT  3.540 1.570 3.780 3.010 ;
        RECT  3.060 1.570 3.780 1.810 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.041  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.610 2.580 17.630 3.020 ;
        RECT  17.310 1.250 17.630 3.020 ;
        RECT  15.750 1.900 17.630 2.140 ;
        RECT  17.230 1.250 17.630 2.140 ;
        RECT  15.300 3.750 17.010 4.150 ;
        RECT  16.610 2.580 17.010 4.150 ;
        RECT  15.750 1.250 16.150 2.140 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.520 1.060 3.020 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.590 2.580 3.300 3.020 ;
        RECT  2.590 2.170 2.830 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.920 5.600 ;
        RECT  17.310 4.410 17.710 5.600 ;
        RECT  16.040 4.620 16.440 5.600 ;
        RECT  14.700 4.590 15.100 5.600 ;
        RECT  13.150 4.620 13.550 5.600 ;
        RECT  10.450 3.960 10.850 5.600 ;
        RECT  9.070 3.960 9.470 5.600 ;
        RECT  5.950 4.240 6.190 5.600 ;
        RECT  5.520 4.240 6.190 4.480 ;
        RECT  4.210 4.620 4.610 5.600 ;
        RECT  1.990 4.620 2.390 5.600 ;
        RECT  0.720 4.560 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.920 0.740 ;
        RECT  16.490 0.000 16.890 1.550 ;
        RECT  15.180 0.000 15.580 0.980 ;
        RECT  13.280 0.000 13.680 1.000 ;
        RECT  9.950 0.000 10.350 1.210 ;
        RECT  5.640 0.000 6.040 0.930 ;
        RECT  4.660 0.000 5.060 0.930 ;
        RECT  0.740 0.000 1.140 1.040 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.340 1.820 ;
        RECT  1.100 1.580 1.340 2.260 ;
        RECT  1.100 2.020 1.790 2.260 ;
        RECT  1.550 2.020 1.790 3.520 ;
        RECT  0.150 3.280 1.790 3.520 ;
        RECT  1.590 1.180 2.350 1.420 ;
        RECT  1.590 1.180 1.830 1.780 ;
        RECT  4.230 2.800 4.480 3.490 ;
        RECT  2.110 3.260 4.350 3.500 ;
        RECT  2.110 1.180 2.350 4.230 ;
        RECT  1.440 3.990 2.350 4.230 ;
        RECT  5.050 1.650 6.030 1.890 ;
        RECT  5.790 2.330 6.440 2.570 ;
        RECT  5.790 1.650 6.030 3.520 ;
        RECT  4.940 3.280 6.030 3.520 ;
        RECT  6.410 1.680 7.040 1.920 ;
        RECT  6.800 1.680 7.040 3.050 ;
        RECT  6.330 2.810 7.040 3.050 ;
        RECT  6.330 2.810 6.570 3.510 ;
        RECT  3.330 1.030 4.260 1.270 ;
        RECT  4.010 1.170 7.530 1.410 ;
        RECT  7.290 1.170 7.530 2.100 ;
        RECT  7.380 1.860 7.620 3.530 ;
        RECT  7.030 3.290 7.620 3.530 ;
        RECT  3.160 3.740 4.740 3.980 ;
        RECT  7.030 3.290 7.270 4.000 ;
        RECT  4.430 3.760 7.270 4.000 ;
        RECT  8.510 1.540 9.090 1.780 ;
        RECT  8.510 1.540 8.750 3.720 ;
        RECT  8.990 3.360 10.150 3.600 ;
        RECT  8.510 3.480 9.230 3.720 ;
        RECT  8.030 0.980 9.710 1.220 ;
        RECT  9.470 0.980 9.710 1.770 ;
        RECT  9.470 1.530 11.130 1.770 ;
        RECT  10.890 1.530 11.130 2.140 ;
        RECT  8.030 0.980 8.270 2.210 ;
        RECT  7.990 1.970 8.230 4.500 ;
        RECT  7.600 4.250 8.230 4.500 ;
        RECT  10.690 0.980 11.610 1.220 ;
        RECT  8.990 2.020 10.550 2.260 ;
        RECT  10.310 2.020 10.550 2.620 ;
        RECT  8.990 2.020 9.230 2.570 ;
        RECT  10.310 2.380 11.610 2.620 ;
        RECT  11.370 0.980 11.610 3.110 ;
        RECT  11.010 2.870 11.610 3.110 ;
        RECT  12.330 1.550 12.910 1.790 ;
        RECT  12.330 1.550 12.570 3.380 ;
        RECT  12.330 2.980 12.780 3.380 ;
        RECT  14.290 2.090 14.530 2.750 ;
        RECT  13.290 2.510 14.530 2.750 ;
        RECT  13.290 2.510 13.530 3.110 ;
        RECT  13.020 2.870 13.530 3.110 ;
        RECT  11.850 1.480 12.090 4.120 ;
        RECT  11.850 3.660 13.260 3.900 ;
        RECT  13.020 2.870 13.260 3.900 ;
        RECT  11.790 3.720 12.190 4.120 ;
        RECT  13.920 0.980 14.880 1.230 ;
        RECT  13.920 0.980 14.160 1.520 ;
        RECT  13.170 1.280 14.160 1.520 ;
        RECT  14.470 0.980 14.880 1.520 ;
        RECT  13.170 1.280 13.410 2.270 ;
        RECT  12.810 2.030 13.410 2.270 ;
        RECT  14.770 1.910 15.450 2.310 ;
        RECT  12.810 2.030 13.050 2.630 ;
        RECT  14.770 1.280 15.010 4.090 ;
        RECT  13.980 3.850 15.010 4.090 ;
        RECT  13.980 3.850 14.220 4.430 ;
    END
END sdcfq4

MACRO sdcfq2
    CLASS CORE ;
    FOREIGN sdcfq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.497  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.020 16.140 2.460 ;
        RECT  15.620 1.990 16.020 2.390 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.122  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 3.700 7.250 4.260 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.338  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.860 3.140 17.300 3.580 ;
        RECT  16.860 1.460 17.130 3.750 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.920 5.600 ;
        RECT  17.450 4.200 17.690 5.600 ;
        RECT  16.150 4.200 16.390 5.600 ;
        RECT  14.830 4.200 15.070 5.600 ;
        RECT  11.810 4.350 12.050 5.600 ;
        RECT  10.450 4.350 10.690 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.920 0.740 ;
        RECT  16.190 0.000 16.590 0.890 ;
        RECT  14.310 0.000 14.710 0.890 ;
        RECT  11.530 0.000 11.770 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.250 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.080 0.570 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.150 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.150 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  10.320 1.750 10.560 3.630 ;
        RECT  10.320 3.130 10.660 3.630 ;
        RECT  10.320 3.390 11.540 3.630 ;
        RECT  9.580 1.270 11.060 1.510 ;
        RECT  10.820 1.270 11.060 2.600 ;
        RECT  10.820 2.360 12.320 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  12.230 1.830 12.810 2.070 ;
        RECT  12.570 1.830 12.810 3.100 ;
        RECT  11.300 2.860 12.810 3.100 ;
        RECT  12.330 2.860 12.570 3.630 ;
        RECT  12.330 3.390 12.900 3.630 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 2.410 8.740 2.810 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 12.530 4.110 ;
        RECT  12.290 3.870 12.530 4.490 ;
        RECT  12.290 4.250 13.150 4.490 ;
        RECT  13.800 1.610 14.050 2.010 ;
        RECT  13.800 1.610 14.040 3.960 ;
        RECT  13.800 3.720 14.380 3.960 ;
        RECT  13.050 1.130 15.000 1.370 ;
        RECT  14.760 1.130 15.000 2.840 ;
        RECT  13.050 1.130 13.290 3.180 ;
        RECT  14.970 2.600 15.370 3.000 ;
        RECT  13.050 2.940 13.560 3.180 ;
        RECT  13.320 2.940 13.560 3.710 ;
        RECT  15.540 1.500 16.620 1.740 ;
        RECT  16.380 1.500 16.620 3.140 ;
        RECT  14.280 2.770 14.520 3.480 ;
        RECT  16.250 2.900 16.490 3.480 ;
        RECT  14.280 3.240 16.490 3.480 ;
        RECT  15.330 3.240 15.730 3.750 ;
    END
END sdcfq2

MACRO sdcfq1
    CLASS CORE ;
    FOREIGN sdcfq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.020 16.140 2.460 ;
        RECT  15.620 1.990 16.020 2.390 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.122  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 3.700 7.250 4.260 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.009  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.860 3.140 17.240 3.750 ;
        RECT  16.860 1.460 17.130 3.750 ;
        END
    END Q
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.360 5.600 ;
        RECT  16.280 4.200 16.520 5.600 ;
        RECT  14.830 4.200 15.070 5.600 ;
        RECT  11.810 4.350 12.050 5.600 ;
        RECT  10.450 4.350 10.690 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.190 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.360 0.740 ;
        RECT  16.270 0.000 16.510 1.190 ;
        RECT  14.310 0.000 14.710 0.890 ;
        RECT  11.530 0.000 11.770 2.050 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.250 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.550 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 2.150 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  8.720 1.730 9.220 2.150 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.980 1.730 9.220 3.450 ;
        RECT  8.860 3.130 9.220 3.450 ;
        RECT  10.320 1.750 10.560 3.630 ;
        RECT  10.320 3.130 10.740 3.630 ;
        RECT  10.320 3.390 11.540 3.630 ;
        RECT  9.580 1.270 11.060 1.510 ;
        RECT  10.820 1.270 11.060 2.600 ;
        RECT  10.820 2.360 12.320 2.600 ;
        RECT  9.580 1.270 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  12.230 1.830 12.810 2.070 ;
        RECT  12.570 1.830 12.810 3.100 ;
        RECT  11.300 2.860 12.810 3.100 ;
        RECT  12.330 2.860 12.570 3.630 ;
        RECT  12.330 3.390 12.900 3.630 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 2.410 8.740 2.810 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 12.530 4.110 ;
        RECT  12.290 3.870 12.530 4.490 ;
        RECT  12.290 4.250 13.150 4.490 ;
        RECT  13.800 1.610 14.050 2.010 ;
        RECT  13.800 1.610 14.040 3.960 ;
        RECT  13.800 3.720 14.380 3.960 ;
        RECT  13.050 1.130 15.000 1.370 ;
        RECT  14.760 1.130 15.000 2.840 ;
        RECT  13.050 1.130 13.290 3.180 ;
        RECT  14.970 2.600 15.370 3.000 ;
        RECT  13.050 2.940 13.560 3.180 ;
        RECT  13.320 2.940 13.560 3.710 ;
        RECT  15.540 1.500 16.620 1.740 ;
        RECT  14.280 2.770 14.520 3.480 ;
        RECT  16.380 1.500 16.620 3.480 ;
        RECT  14.280 3.240 16.620 3.480 ;
        RECT  15.460 3.240 15.860 3.750 ;
    END
END sdcfq1

MACRO sdcfb4
    CLASS CORE ;
    FOREIGN sdcfb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.377  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.580 7.510 3.020 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.459  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.180 2.590 15.710 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.453  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.600 2.820 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.771  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.960 3.750 14.620 3.990 ;
        RECT  12.800 1.630 14.590 1.870 ;
        RECT  13.960 1.630 14.200 3.990 ;
        RECT  12.870 3.270 14.200 3.640 ;
        RECT  12.800 1.630 14.200 1.890 ;
        RECT  12.870 3.270 13.270 3.840 ;
        RECT  12.380 3.270 14.200 3.580 ;
        RECT  12.380 3.140 12.840 3.580 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.669  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.580 3.840 19.320 4.080 ;
        RECT  17.140 1.820 19.020 2.060 ;
        RECT  18.620 1.560 19.020 2.060 ;
        RECT  17.980 2.580 18.420 3.020 ;
        RECT  18.090 1.820 18.330 4.080 ;
        RECT  17.140 1.560 17.540 2.060 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.670 3.070 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.210 3.020 ;
        RECT  3.970 2.210 4.210 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.160 5.600 ;
        RECT  19.650 3.080 19.890 5.600 ;
        RECT  18.360 4.560 18.760 5.600 ;
        RECT  16.960 4.590 17.360 5.600 ;
        RECT  15.020 4.710 15.420 5.600 ;
        RECT  13.660 4.710 14.060 5.600 ;
        RECT  12.300 4.710 12.700 5.600 ;
        RECT  10.900 4.710 11.300 5.600 ;
        RECT  7.920 4.710 8.320 5.600 ;
        RECT  6.740 4.710 7.130 5.600 ;
        RECT  3.260 4.520 3.660 5.600 ;
        RECT  0.780 4.620 1.180 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.160 0.740 ;
        RECT  19.440 0.000 19.680 1.420 ;
        RECT  17.960 0.000 18.200 1.420 ;
        RECT  15.480 0.000 15.880 0.890 ;
        RECT  13.540 0.000 13.940 0.890 ;
        RECT  7.290 0.000 7.530 1.650 ;
        RECT  3.180 1.070 3.780 1.320 ;
        RECT  3.540 0.000 3.780 1.320 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.340 1.820 ;
        RECT  1.100 1.580 1.340 2.910 ;
        RECT  1.000 2.700 1.240 3.590 ;
        RECT  0.150 3.350 1.240 3.590 ;
        RECT  1.590 2.100 3.510 2.340 ;
        RECT  1.590 1.760 1.830 3.230 ;
        RECT  1.530 3.070 1.770 3.670 ;
        RECT  1.980 0.980 2.770 1.220 ;
        RECT  2.530 0.980 2.770 1.860 ;
        RECT  2.530 1.620 4.700 1.860 ;
        RECT  4.460 1.070 4.700 3.650 ;
        RECT  2.150 3.330 4.790 3.570 ;
        RECT  4.460 3.250 4.790 3.650 ;
        RECT  4.410 3.330 4.790 3.650 ;
        RECT  5.710 1.500 6.290 1.740 ;
        RECT  5.710 1.500 5.950 2.270 ;
        RECT  5.700 2.190 5.940 3.510 ;
        RECT  5.700 3.270 7.730 3.510 ;
        RECT  5.220 1.420 5.470 1.740 ;
        RECT  5.220 1.420 5.460 4.140 ;
        RECT  5.220 3.750 8.210 3.990 ;
        RECT  7.970 2.630 8.210 3.990 ;
        RECT  5.150 3.790 5.540 4.140 ;
        RECT  6.240 2.060 8.300 2.300 ;
        RECT  8.060 1.440 8.300 2.300 ;
        RECT  8.090 2.150 8.750 2.390 ;
        RECT  6.240 2.060 6.480 2.630 ;
        RECT  8.510 2.150 8.750 3.090 ;
        RECT  8.510 2.850 9.010 3.090 ;
        RECT  8.770 2.850 9.010 3.740 ;
        RECT  9.480 1.530 10.070 1.770 ;
        RECT  9.830 1.530 10.070 3.370 ;
        RECT  9.830 3.130 10.570 3.370 ;
        RECT  8.740 1.470 9.230 1.870 ;
        RECT  11.000 2.080 11.960 2.320 ;
        RECT  8.990 1.470 9.230 2.610 ;
        RECT  8.990 2.370 9.490 2.610 ;
        RECT  9.250 2.370 9.490 3.990 ;
        RECT  11.000 2.080 11.240 3.990 ;
        RECT  9.250 3.750 11.240 3.990 ;
        RECT  10.310 1.520 12.440 1.760 ;
        RECT  12.200 2.240 13.310 2.480 ;
        RECT  12.200 1.520 12.440 2.810 ;
        RECT  11.790 2.570 12.440 2.810 ;
        RECT  10.310 1.520 10.550 2.870 ;
        RECT  11.790 2.570 12.030 3.980 ;
        RECT  11.530 3.580 12.030 3.980 ;
        RECT  8.500 0.980 13.300 1.220 ;
        RECT  13.070 1.130 15.210 1.370 ;
        RECT  14.970 1.130 15.210 2.350 ;
        RECT  14.700 2.110 16.080 2.350 ;
        RECT  15.900 2.180 16.400 2.420 ;
        RECT  14.700 2.110 14.940 3.520 ;
        RECT  14.700 3.280 15.930 3.520 ;
        RECT  15.690 3.280 15.930 3.970 ;
        RECT  16.610 0.980 17.190 1.220 ;
        RECT  16.250 1.640 16.850 1.880 ;
        RECT  16.610 0.980 16.850 1.880 ;
        RECT  16.640 1.710 16.880 2.970 ;
        RECT  16.400 2.730 16.640 4.460 ;
        RECT  5.970 4.230 8.890 4.470 ;
        RECT  9.710 4.230 16.640 4.460 ;
        RECT  5.490 4.380 16.630 4.470 ;
        RECT  5.490 4.380 6.240 4.620 ;
        RECT  8.620 4.380 10.000 4.620 ;
    END
END sdcfb4

MACRO sdcfb2
    CLASS CORE ;
    FOREIGN sdcfb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.395  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.580 7.510 3.020 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.456  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.810 2.020 14.500 2.460 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.453  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.600 2.820 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.343  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.140 1.610 13.380 3.380 ;
        RECT  12.730 3.140 13.270 3.840 ;
        RECT  12.800 1.610 13.380 1.850 ;
        RECT  12.380 3.140 13.270 3.580 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.585  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.230 2.520 17.130 3.160 ;
        RECT  16.890 1.420 17.130 3.160 ;
        RECT  16.230 2.520 16.630 3.550 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.670 3.070 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.210 3.020 ;
        RECT  3.970 2.210 4.210 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.360 5.600 ;
        RECT  16.890 3.820 17.130 5.600 ;
        RECT  15.570 3.990 15.810 5.600 ;
        RECT  13.600 4.710 14.000 5.600 ;
        RECT  12.240 4.710 12.640 5.600 ;
        RECT  10.840 4.710 11.240 5.600 ;
        RECT  7.920 4.710 8.320 5.600 ;
        RECT  6.740 4.710 7.130 5.600 ;
        RECT  3.260 4.520 3.660 5.600 ;
        RECT  0.780 4.620 1.180 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.360 0.740 ;
        RECT  16.050 0.000 16.450 0.980 ;
        RECT  13.130 0.000 13.530 0.890 ;
        RECT  7.210 0.000 7.610 1.650 ;
        RECT  3.180 1.070 3.870 1.320 ;
        RECT  3.610 0.000 3.870 1.320 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.340 1.820 ;
        RECT  1.100 1.580 1.340 2.910 ;
        RECT  1.000 2.700 1.240 3.590 ;
        RECT  0.150 3.350 1.240 3.590 ;
        RECT  1.590 2.100 3.510 2.340 ;
        RECT  1.590 1.760 1.830 3.230 ;
        RECT  1.530 3.070 1.770 3.670 ;
        RECT  1.980 0.980 2.770 1.220 ;
        RECT  2.530 0.980 2.770 1.860 ;
        RECT  2.530 1.620 4.700 1.860 ;
        RECT  4.460 1.070 4.700 3.570 ;
        RECT  4.390 3.250 4.800 3.570 ;
        RECT  4.460 3.180 4.800 3.570 ;
        RECT  2.150 3.330 4.800 3.570 ;
        RECT  5.710 1.500 6.290 1.740 ;
        RECT  5.710 1.500 5.950 2.270 ;
        RECT  5.700 2.190 5.940 3.510 ;
        RECT  5.700 3.270 7.730 3.510 ;
        RECT  5.220 1.420 5.470 1.740 ;
        RECT  5.220 1.420 5.460 4.140 ;
        RECT  5.220 3.750 8.210 3.990 ;
        RECT  7.970 2.630 8.210 3.990 ;
        RECT  5.140 3.770 5.540 4.140 ;
        RECT  8.060 1.440 8.300 2.340 ;
        RECT  6.240 2.100 8.690 2.340 ;
        RECT  6.240 2.100 6.480 2.670 ;
        RECT  8.450 2.100 8.690 3.090 ;
        RECT  8.450 2.850 8.950 3.090 ;
        RECT  8.710 2.850 8.950 3.740 ;
        RECT  9.480 1.510 10.070 1.780 ;
        RECT  9.830 1.510 10.070 3.370 ;
        RECT  9.830 3.130 10.500 3.370 ;
        RECT  8.740 1.460 9.230 1.860 ;
        RECT  10.950 2.120 11.980 2.360 ;
        RECT  8.990 1.460 9.230 2.610 ;
        RECT  8.990 2.370 9.590 2.610 ;
        RECT  9.350 2.370 9.590 4.070 ;
        RECT  9.350 3.670 9.710 4.070 ;
        RECT  10.950 2.120 11.190 3.990 ;
        RECT  9.350 3.750 11.190 3.990 ;
        RECT  9.350 3.750 9.760 4.070 ;
        RECT  10.310 1.520 12.460 1.760 ;
        RECT  12.220 2.240 12.770 2.480 ;
        RECT  10.310 1.520 10.550 2.870 ;
        RECT  12.220 1.520 12.460 2.900 ;
        RECT  11.790 2.660 12.460 2.900 ;
        RECT  11.790 2.660 12.030 3.980 ;
        RECT  11.470 3.570 12.030 3.980 ;
        RECT  8.500 0.980 12.890 1.220 ;
        RECT  12.660 1.130 14.030 1.370 ;
        RECT  13.780 1.130 14.030 1.770 ;
        RECT  13.780 1.530 14.950 1.770 ;
        RECT  14.760 1.620 15.240 1.860 ;
        RECT  14.990 1.620 15.240 2.940 ;
        RECT  14.290 2.700 15.240 2.940 ;
        RECT  14.290 2.700 14.530 3.800 ;
        RECT  14.660 0.980 15.720 1.220 ;
        RECT  15.250 0.980 15.720 1.380 ;
        RECT  15.480 0.980 15.720 3.550 ;
        RECT  14.920 3.310 15.720 3.550 ;
        RECT  14.920 3.310 15.320 3.650 ;
        RECT  12.670 4.080 15.240 4.320 ;
        RECT  15.000 3.310 15.240 4.320 ;
        RECT  5.970 4.230 8.890 4.470 ;
        RECT  10.150 4.230 12.940 4.470 ;
        RECT  5.490 4.380 6.240 4.620 ;
        RECT  8.620 4.380 10.410 4.620 ;
    END
END sdcfb2

MACRO sdcfb1
    CLASS CORE ;
    FOREIGN sdcfb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.458  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.100 2.480 15.620 3.020 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.395  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.580 7.510 3.020 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.453  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.600 2.820 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.127  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.730 3.720 13.290 3.960 ;
        RECT  12.380 3.140 13.280 3.380 ;
        RECT  13.040 1.520 13.280 3.380 ;
        RECT  12.870 1.520 13.280 1.920 ;
        RECT  12.730 3.140 12.970 3.960 ;
        RECT  12.380 3.140 12.970 3.580 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.300 2.580 16.680 3.020 ;
        RECT  16.330 1.700 16.570 4.110 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.670 3.070 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.210 3.020 ;
        RECT  3.970 2.210 4.210 3.020 ;
        END
    END SD
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  15.680 4.480 16.080 5.600 ;
        RECT  14.170 4.400 14.570 5.600 ;
        RECT  12.300 4.710 12.700 5.600 ;
        RECT  10.900 4.710 11.300 5.600 ;
        RECT  7.920 4.710 8.320 5.600 ;
        RECT  6.740 4.710 7.130 5.600 ;
        RECT  3.260 4.520 3.660 5.600 ;
        RECT  0.780 4.620 1.180 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  15.900 0.000 16.300 0.890 ;
        RECT  14.220 0.000 14.620 0.890 ;
        RECT  10.380 0.000 10.760 0.890 ;
        RECT  10.350 0.000 10.760 0.870 ;
        RECT  7.210 0.000 7.610 1.650 ;
        RECT  3.180 1.080 3.770 1.320 ;
        RECT  3.530 0.000 3.770 1.320 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.340 1.820 ;
        RECT  1.100 1.580 1.340 2.910 ;
        RECT  1.000 2.700 1.240 3.590 ;
        RECT  0.150 3.350 1.240 3.590 ;
        RECT  1.590 2.100 3.510 2.340 ;
        RECT  1.590 1.680 1.830 3.230 ;
        RECT  1.530 3.070 1.770 3.670 ;
        RECT  1.980 0.980 2.770 1.220 ;
        RECT  2.530 0.980 2.770 1.860 ;
        RECT  2.530 1.620 4.700 1.860 ;
        RECT  4.460 1.070 4.700 3.670 ;
        RECT  2.150 3.330 4.790 3.570 ;
        RECT  4.460 3.240 4.790 3.670 ;
        RECT  4.390 3.330 4.790 3.670 ;
        RECT  5.710 1.500 6.290 1.740 ;
        RECT  5.710 1.500 5.950 2.270 ;
        RECT  5.700 2.190 5.940 3.510 ;
        RECT  5.700 3.270 7.730 3.510 ;
        RECT  5.230 1.420 5.470 1.970 ;
        RECT  5.220 1.770 5.460 4.140 ;
        RECT  7.970 2.630 8.210 3.990 ;
        RECT  5.140 3.750 8.210 3.990 ;
        RECT  5.140 3.750 5.540 4.140 ;
        RECT  6.240 2.060 8.300 2.300 ;
        RECT  8.060 1.440 8.300 2.300 ;
        RECT  8.090 2.150 8.750 2.390 ;
        RECT  6.240 2.060 6.480 2.660 ;
        RECT  8.510 2.150 8.750 3.350 ;
        RECT  8.510 3.110 9.010 3.350 ;
        RECT  8.770 3.110 9.010 3.740 ;
        RECT  9.560 1.470 9.800 2.390 ;
        RECT  9.560 2.150 10.070 2.390 ;
        RECT  9.830 2.150 10.070 3.370 ;
        RECT  9.830 3.130 10.570 3.370 ;
        RECT  8.740 1.470 9.230 1.870 ;
        RECT  11.070 2.130 12.020 2.370 ;
        RECT  8.990 1.470 9.230 2.870 ;
        RECT  8.990 2.630 9.590 2.870 ;
        RECT  11.070 2.130 11.310 3.450 ;
        RECT  9.350 2.630 9.590 4.070 ;
        RECT  11.000 3.220 11.240 3.990 ;
        RECT  9.350 3.670 11.240 3.990 ;
        RECT  9.350 3.670 9.770 4.070 ;
        RECT  11.450 1.520 12.140 1.790 ;
        RECT  10.310 1.650 11.650 1.890 ;
        RECT  11.930 1.640 12.500 1.890 ;
        RECT  12.260 2.160 12.800 2.560 ;
        RECT  12.260 1.640 12.500 2.850 ;
        RECT  11.870 2.610 12.500 2.850 ;
        RECT  10.310 1.650 10.550 2.870 ;
        RECT  11.870 2.610 12.110 3.990 ;
        RECT  11.530 3.730 12.110 3.990 ;
        RECT  8.500 1.030 10.160 1.220 ;
        RECT  8.500 1.060 10.180 1.220 ;
        RECT  8.500 1.080 10.220 1.220 ;
        RECT  10.990 1.040 13.980 1.240 ;
        RECT  8.500 0.980 10.130 1.220 ;
        RECT  11.950 1.000 13.980 1.240 ;
        RECT  9.980 1.130 12.330 1.280 ;
        RECT  9.980 1.130 11.230 1.310 ;
        RECT  10.040 1.130 11.230 1.410 ;
        RECT  14.700 1.720 15.350 2.230 ;
        RECT  14.200 2.090 14.910 2.330 ;
        RECT  14.200 2.090 14.440 3.550 ;
        RECT  14.200 3.310 15.020 3.550 ;
        RECT  14.780 3.310 15.020 4.230 ;
        RECT  14.780 3.990 15.380 4.230 ;
        RECT  14.910 0.980 15.540 1.230 ;
        RECT  14.910 0.980 15.150 1.480 ;
        RECT  14.220 1.240 15.150 1.480 ;
        RECT  14.220 1.240 14.460 1.750 ;
        RECT  13.580 1.510 14.460 1.750 ;
        RECT  13.580 1.510 13.980 1.850 ;
        RECT  5.970 4.230 8.890 4.470 ;
        RECT  10.100 4.230 13.920 4.470 ;
        RECT  13.660 1.510 13.920 4.470 ;
        RECT  5.490 4.380 6.240 4.620 ;
        RECT  8.620 4.380 10.390 4.620 ;
    END
END sdcfb1

MACRO sdbrb4
    CLASS CORE ;
    FOREIGN sdbrb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.406  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.750 2.020 13.380 2.760 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.456  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  21.340 3.140 21.780 3.580 ;
        RECT  21.540 2.560 21.780 3.580 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.870 1.960 4.110 2.530 ;
        RECT  3.420 2.580 3.920 3.020 ;
        RECT  3.660 2.290 3.920 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.638  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.180 3.550 17.140 3.790 ;
        RECT  16.850 1.880 17.140 3.790 ;
        RECT  16.140 2.580 17.140 3.020 ;
        RECT  16.720 1.880 17.140 3.020 ;
        RECT  14.750 1.880 17.140 2.120 ;
        RECT  16.230 1.560 16.470 2.120 ;
        RECT  14.750 1.310 14.990 2.120 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.787  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.240 1.540 19.480 4.060 ;
        RECT  17.710 1.530 19.430 1.770 ;
        RECT  17.920 2.340 19.480 2.580 ;
        RECT  19.190 1.050 19.430 2.580 ;
        RECT  18.540 1.540 19.480 2.580 ;
        RECT  17.920 2.340 18.160 4.060 ;
        RECT  17.710 1.100 17.950 1.770 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.370 2.180 3.020 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.940 2.680 8.380 3.080 ;
        RECT  7.340 2.580 7.950 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 22.400 5.600 ;
        RECT  21.120 4.400 21.520 5.600 ;
        RECT  19.790 2.850 20.030 5.600 ;
        RECT  18.480 2.980 18.720 5.600 ;
        RECT  17.120 4.520 17.520 5.600 ;
        RECT  15.760 4.520 16.160 5.600 ;
        RECT  14.400 4.710 14.800 5.600 ;
        RECT  13.180 4.710 13.580 5.600 ;
        RECT  11.350 4.710 11.750 5.600 ;
        RECT  8.680 4.710 9.080 5.600 ;
        RECT  6.420 4.710 6.820 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.720 3.550 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 22.400 0.740 ;
        RECT  20.550 0.000 20.970 1.220 ;
        RECT  18.370 0.000 18.770 1.290 ;
        RECT  16.890 0.000 17.290 1.620 ;
        RECT  15.410 0.000 15.810 1.640 ;
        RECT  13.900 0.000 14.300 1.260 ;
        RECT  11.880 0.000 12.280 1.260 ;
        RECT  9.750 0.000 10.150 0.820 ;
        RECT  7.420 0.000 7.660 1.720 ;
        RECT  3.320 0.000 3.560 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.430 1.270 1.670 ;
        RECT  1.030 1.430 1.270 3.310 ;
        RECT  1.030 2.520 1.450 2.940 ;
        RECT  1.030 2.520 1.290 3.310 ;
        RECT  0.230 3.070 1.290 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.510 1.700 2.600 1.940 ;
        RECT  2.360 1.920 3.400 2.160 ;
        RECT  2.420 1.920 2.660 3.460 ;
        RECT  1.540 3.260 2.570 3.500 ;
        RECT  1.540 3.260 1.780 4.000 ;
        RECT  2.040 1.010 3.080 1.250 ;
        RECT  2.840 1.010 3.080 1.680 ;
        RECT  4.520 1.050 4.760 1.600 ;
        RECT  2.840 1.440 4.750 1.680 ;
        RECT  4.520 1.050 4.590 3.010 ;
        RECT  4.350 1.440 4.530 3.940 ;
        RECT  4.290 2.770 4.530 3.940 ;
        RECT  2.710 3.700 4.530 3.940 ;
        RECT  2.710 3.700 2.950 4.620 ;
        RECT  1.990 4.380 2.950 4.620 ;
        RECT  4.990 1.670 5.230 2.230 ;
        RECT  4.830 1.990 5.070 3.390 ;
        RECT  4.770 3.200 5.010 4.620 ;
        RECT  4.770 4.380 5.770 4.620 ;
        RECT  5.950 1.460 6.540 1.700 ;
        RECT  5.790 3.010 6.190 3.410 ;
        RECT  5.950 1.460 6.190 4.060 ;
        RECT  5.940 3.740 6.190 4.060 ;
        RECT  5.940 3.820 7.590 4.060 ;
        RECT  5.270 0.980 7.020 1.220 ;
        RECT  5.270 0.980 5.710 1.380 ;
        RECT  6.780 0.980 7.020 2.200 ;
        RECT  6.780 1.960 8.620 2.200 ;
        RECT  8.380 2.200 8.860 2.440 ;
        RECT  5.470 0.980 5.710 2.710 ;
        RECT  8.620 2.200 8.860 2.990 ;
        RECT  8.620 2.750 9.240 2.990 ;
        RECT  5.310 2.470 5.550 3.810 ;
        RECT  5.250 3.580 5.490 4.140 ;
        RECT  9.010 1.580 9.410 1.990 ;
        RECT  9.160 1.580 9.410 2.510 ;
        RECT  9.160 2.270 9.720 2.510 ;
        RECT  6.430 2.440 6.670 3.570 ;
        RECT  6.430 3.330 9.720 3.570 ;
        RECT  9.480 2.270 9.720 3.650 ;
        RECT  9.260 3.250 9.720 3.650 ;
        RECT  7.900 1.100 11.410 1.340 ;
        RECT  7.900 1.020 8.320 1.430 ;
        RECT  11.170 1.100 11.410 1.740 ;
        RECT  11.170 1.500 11.950 1.740 ;
        RECT  11.710 1.500 11.950 2.200 ;
        RECT  10.440 1.650 10.890 2.050 ;
        RECT  10.440 2.930 10.850 3.330 ;
        RECT  10.440 1.650 10.680 3.330 ;
        RECT  10.610 3.260 12.280 3.500 ;
        RECT  8.050 4.230 9.560 4.470 ;
        RECT  10.880 4.230 12.210 4.470 ;
        RECT  7.550 4.350 8.290 4.590 ;
        RECT  9.320 4.380 11.120 4.620 ;
        RECT  11.980 4.380 12.810 4.620 ;
        RECT  13.280 0.980 13.520 1.780 ;
        RECT  12.270 1.540 14.200 1.780 ;
        RECT  13.960 2.360 15.900 2.600 ;
        RECT  10.950 2.290 11.370 2.690 ;
        RECT  11.130 2.290 11.370 2.950 ;
        RECT  12.270 1.540 12.510 2.950 ;
        RECT  11.130 2.710 12.510 2.950 ;
        RECT  13.960 1.540 14.200 3.450 ;
        RECT  12.580 3.210 14.200 3.450 ;
        RECT  9.750 1.630 10.200 2.030 ;
        RECT  9.960 1.630 10.200 4.140 ;
        RECT  9.960 3.740 13.420 3.990 ;
        RECT  13.180 3.740 13.420 4.270 ;
        RECT  9.960 3.740 10.380 4.140 ;
        RECT  17.440 2.010 17.680 4.270 ;
        RECT  13.180 4.030 17.680 4.270 ;
        RECT  19.720 1.010 20.210 1.410 ;
        RECT  19.720 1.010 19.960 2.610 ;
        RECT  19.720 2.370 20.580 2.610 ;
        RECT  20.340 2.370 20.580 3.410 ;
        RECT  20.340 3.170 20.930 3.410 ;
        RECT  21.290 1.330 22.260 1.570 ;
        RECT  20.210 1.890 22.260 2.130 ;
        RECT  21.860 3.810 22.260 4.210 ;
        RECT  22.020 1.330 22.260 4.210 ;
        RECT  21.850 3.820 22.260 4.210 ;
    END
END sdbrb4

MACRO sdbrb2
    CLASS CORE ;
    FOREIGN sdbrb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.420 2.340 17.860 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.197  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  20.550 1.650 20.790 3.100 ;
        RECT  20.220 2.860 20.660 3.580 ;
        RECT  20.060 1.650 20.790 1.890 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.196  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.720 3.130 19.250 3.450 ;
        RECT  18.720 1.570 18.980 3.450 ;
        RECT  18.540 2.580 18.980 3.020 ;
        RECT  18.680 1.570 18.980 3.020 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.257  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.331  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.380 2.020 12.880 2.520 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 21.280 5.600 ;
        RECT  20.810 4.170 21.050 5.600 ;
        RECT  19.500 4.170 19.740 5.600 ;
        RECT  18.190 4.170 18.430 5.600 ;
        RECT  16.890 4.150 17.130 5.600 ;
        RECT  15.500 3.920 15.740 5.600 ;
        RECT  12.700 4.350 12.940 5.600 ;
        RECT  11.810 4.400 12.050 5.600 ;
        RECT  10.450 4.400 10.690 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.530 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 21.280 0.740 ;
        RECT  20.810 0.000 21.050 1.400 ;
        RECT  19.390 0.000 19.630 1.400 ;
        RECT  18.010 0.000 18.250 1.140 ;
        RECT  15.990 0.000 16.390 0.890 ;
        RECT  11.530 0.000 11.770 1.890 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.550 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 1.980 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.940 1.580 9.180 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.480 4.110 ;
        RECT  10.330 1.590 10.570 3.630 ;
        RECT  10.330 3.130 10.740 3.630 ;
        RECT  10.330 3.390 11.540 3.630 ;
        RECT  9.580 1.110 11.060 1.350 ;
        RECT  10.820 1.110 11.060 2.440 ;
        RECT  10.820 2.200 12.140 2.440 ;
        RECT  9.580 1.110 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  12.730 1.520 13.360 1.760 ;
        RECT  11.300 2.860 12.020 3.100 ;
        RECT  11.780 2.860 12.020 3.400 ;
        RECT  13.120 1.520 13.360 3.400 ;
        RECT  11.780 3.160 13.640 3.400 ;
        RECT  13.240 3.140 13.640 3.480 ;
        RECT  9.850 3.870 13.690 4.110 ;
        RECT  13.450 3.870 13.690 4.500 ;
        RECT  13.450 4.260 14.160 4.500 ;
        RECT  14.440 1.670 15.000 1.910 ;
        RECT  14.760 1.670 15.000 3.710 ;
        RECT  14.760 3.390 16.460 3.630 ;
        RECT  14.760 3.390 15.160 3.710 ;
        RECT  13.760 1.130 16.510 1.370 ;
        RECT  16.270 1.130 16.510 2.520 ;
        RECT  16.270 2.120 16.670 2.520 ;
        RECT  13.760 1.130 14.000 2.900 ;
        RECT  13.760 2.660 14.330 2.900 ;
        RECT  14.090 2.660 14.330 3.710 ;
        RECT  16.940 1.500 17.620 1.740 ;
        RECT  19.560 2.180 20.310 2.420 ;
        RECT  15.650 2.250 15.890 3.020 ;
        RECT  15.650 2.780 17.180 3.020 ;
        RECT  16.940 1.500 17.180 3.630 ;
        RECT  16.940 3.390 18.300 3.630 ;
        RECT  18.060 3.390 18.300 3.930 ;
        RECT  19.560 2.180 19.800 3.930 ;
        RECT  18.060 3.690 19.800 3.930 ;
    END
END sdbrb2

MACRO sdbrb1
    CLASS CORE ;
    FOREIGN sdbrb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.420 2.340 17.860 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.840 3.700 7.250 4.550 ;
        RECT  6.780 3.700 7.250 4.200 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.370 4.380 3.660 4.620 ;
        RECT  3.420 3.700 3.660 4.620 ;
        RECT  2.030 4.170 2.610 4.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.264  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  20.040 3.390 20.550 3.710 ;
        RECT  20.040 1.290 20.400 3.710 ;
        RECT  19.620 1.290 20.400 1.900 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.122  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.440 3.390 19.280 3.630 ;
        RECT  18.440 3.140 18.980 3.630 ;
        RECT  18.440 1.210 18.720 3.630 ;
        RECT  18.130 1.210 18.720 1.530 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.257  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.640 1.060 3.160 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.700 5.540 4.140 ;
        RECT  4.860 4.210 5.240 4.610 ;
        RECT  5.000 3.900 5.240 4.610 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.331  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.380 2.020 12.880 2.520 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.720 5.600 ;
        RECT  19.490 4.390 19.730 5.600 ;
        RECT  18.220 4.390 18.460 5.600 ;
        RECT  16.890 4.150 17.130 5.600 ;
        RECT  15.500 3.920 15.740 5.600 ;
        RECT  12.700 4.350 12.940 5.600 ;
        RECT  11.810 4.400 12.050 5.600 ;
        RECT  10.450 4.400 10.690 5.600 ;
        RECT  7.490 3.310 7.730 5.600 ;
        RECT  6.300 4.390 6.540 5.600 ;
        RECT  4.610 3.120 4.850 3.700 ;
        RECT  4.380 3.460 4.620 5.600 ;
        RECT  1.710 4.710 2.090 5.600 ;
        RECT  0.970 4.530 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.720 0.740 ;
        RECT  18.880 0.000 19.280 1.030 ;
        RECT  15.990 0.000 16.390 0.890 ;
        RECT  11.530 0.000 11.770 1.890 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  4.560 0.000 4.960 0.890 ;
        RECT  1.800 0.000 2.040 1.200 ;
        RECT  0.970 0.000 1.210 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.980 0.710 1.220 ;
        RECT  0.470 0.980 0.710 2.400 ;
        RECT  0.140 2.160 1.640 2.400 ;
        RECT  1.320 2.160 1.640 2.550 ;
        RECT  0.140 2.160 0.380 4.490 ;
        RECT  0.140 4.170 0.550 4.490 ;
        RECT  2.360 1.610 2.630 2.010 ;
        RECT  2.360 1.610 2.600 3.450 ;
        RECT  0.950 1.680 2.120 1.920 ;
        RECT  1.880 1.680 2.120 3.930 ;
        RECT  0.920 3.460 2.120 3.700 ;
        RECT  1.880 3.690 3.170 3.930 ;
        RECT  2.850 3.690 3.170 4.140 ;
        RECT  3.710 1.610 4.190 1.930 ;
        RECT  3.710 1.610 3.950 3.130 ;
        RECT  3.840 2.890 4.080 3.450 ;
        RECT  5.090 1.610 5.550 1.940 ;
        RECT  4.190 2.380 5.330 2.620 ;
        RECT  5.090 1.610 5.330 3.340 ;
        RECT  5.090 3.100 5.670 3.340 ;
        RECT  5.570 2.370 6.170 2.610 ;
        RECT  5.930 1.630 6.170 3.940 ;
        RECT  5.820 3.700 6.060 4.620 ;
        RECT  5.480 4.380 6.060 4.620 ;
        RECT  6.740 2.380 7.990 2.620 ;
        RECT  6.740 1.770 6.980 3.450 ;
        RECT  3.100 1.130 8.960 1.370 ;
        RECT  8.720 1.130 8.960 1.980 ;
        RECT  3.100 1.130 3.370 2.000 ;
        RECT  3.100 1.130 3.340 3.450 ;
        RECT  8.940 1.580 9.180 3.450 ;
        RECT  8.020 1.770 8.470 2.090 ;
        RECT  8.230 1.770 8.470 4.110 ;
        RECT  8.230 3.870 9.480 4.110 ;
        RECT  10.330 1.590 10.570 3.630 ;
        RECT  10.330 3.130 10.740 3.630 ;
        RECT  10.330 3.390 11.540 3.630 ;
        RECT  9.580 1.110 11.060 1.350 ;
        RECT  10.820 1.110 11.060 2.440 ;
        RECT  10.820 2.200 12.140 2.440 ;
        RECT  9.580 1.110 9.820 3.450 ;
        RECT  9.580 3.130 10.000 3.450 ;
        RECT  12.730 1.520 13.360 1.760 ;
        RECT  11.300 2.860 12.020 3.100 ;
        RECT  11.780 2.860 12.020 3.400 ;
        RECT  13.120 1.520 13.360 3.400 ;
        RECT  11.780 3.160 13.640 3.400 ;
        RECT  13.240 3.140 13.640 3.480 ;
        RECT  9.850 3.870 13.690 4.110 ;
        RECT  13.450 3.870 13.690 4.500 ;
        RECT  13.450 4.260 14.160 4.500 ;
        RECT  14.440 1.670 15.000 1.910 ;
        RECT  14.760 1.670 15.000 3.710 ;
        RECT  14.760 3.390 16.460 3.630 ;
        RECT  14.760 3.390 15.160 3.710 ;
        RECT  13.760 1.130 16.510 1.370 ;
        RECT  16.270 1.130 16.510 2.520 ;
        RECT  16.270 2.120 16.670 2.520 ;
        RECT  13.760 1.130 14.000 2.900 ;
        RECT  13.760 2.660 14.330 2.900 ;
        RECT  14.090 2.660 14.330 3.710 ;
        RECT  16.940 1.500 17.620 1.740 ;
        RECT  15.650 2.250 15.890 3.020 ;
        RECT  15.650 2.780 17.180 3.020 ;
        RECT  16.940 1.500 17.180 3.630 ;
        RECT  16.940 3.390 18.130 3.630 ;
        RECT  17.880 3.390 18.130 4.120 ;
        RECT  19.520 2.710 19.760 4.120 ;
        RECT  17.880 3.880 19.760 4.120 ;
    END
END sdbrb1

MACRO sdbfb4
    CLASS CORE ;
    FOREIGN sdbfb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.406  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.750 2.020 13.380 2.760 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.456  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  21.230 3.140 21.780 3.580 ;
        RECT  21.370 2.560 21.770 3.580 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.870 1.960 4.110 2.530 ;
        RECT  3.420 2.580 3.920 3.020 ;
        RECT  3.660 2.290 3.920 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.621  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.180 3.550 17.200 3.790 ;
        RECT  16.860 1.880 17.200 3.790 ;
        RECT  16.140 2.580 17.200 3.020 ;
        RECT  16.850 1.880 17.200 3.020 ;
        RECT  14.750 1.880 17.200 2.120 ;
        RECT  16.230 1.260 16.470 2.120 ;
        RECT  14.750 1.310 14.990 2.120 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.733  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.240 2.500 19.480 4.060 ;
        RECT  17.710 1.530 19.430 1.770 ;
        RECT  19.190 1.100 19.430 1.770 ;
        RECT  17.920 2.500 19.480 2.740 ;
        RECT  18.540 1.530 18.980 2.740 ;
        RECT  17.920 2.500 18.160 4.060 ;
        RECT  17.710 1.100 17.950 1.770 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.730 2.370 2.180 3.020 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.940 2.680 8.360 3.080 ;
        RECT  7.340 2.580 7.950 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 22.400 5.600 ;
        RECT  21.000 4.400 21.400 5.600 ;
        RECT  19.790 2.850 20.030 5.600 ;
        RECT  18.480 2.980 18.720 5.600 ;
        RECT  17.120 4.520 17.520 5.600 ;
        RECT  15.760 4.520 16.160 5.600 ;
        RECT  14.400 4.710 14.800 5.600 ;
        RECT  13.180 4.710 13.580 5.600 ;
        RECT  11.350 4.710 11.750 5.600 ;
        RECT  8.680 4.710 9.080 5.600 ;
        RECT  6.420 4.710 6.820 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.720 3.550 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 22.400 0.740 ;
        RECT  20.650 0.000 21.050 1.220 ;
        RECT  18.370 0.000 18.770 1.290 ;
        RECT  16.890 0.000 17.290 1.620 ;
        RECT  15.410 0.000 15.810 1.640 ;
        RECT  13.900 0.000 14.300 1.260 ;
        RECT  11.960 0.000 12.200 1.260 ;
        RECT  9.800 0.000 10.200 0.820 ;
        RECT  7.420 0.000 7.660 1.720 ;
        RECT  3.320 0.000 3.560 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.430 1.120 1.670 ;
        RECT  0.880 1.430 1.120 2.520 ;
        RECT  1.050 2.280 1.350 2.940 ;
        RECT  1.050 2.530 1.450 2.940 ;
        RECT  1.050 2.280 1.290 3.310 ;
        RECT  0.230 3.070 1.290 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.510 1.700 2.600 1.940 ;
        RECT  2.360 1.920 3.400 2.160 ;
        RECT  2.420 1.920 2.660 3.460 ;
        RECT  1.540 3.260 2.570 3.500 ;
        RECT  1.540 3.260 1.780 4.000 ;
        RECT  2.040 1.010 3.080 1.250 ;
        RECT  2.840 1.010 3.080 1.680 ;
        RECT  4.520 1.080 4.760 1.600 ;
        RECT  2.840 1.440 4.750 1.680 ;
        RECT  4.520 1.080 4.590 3.010 ;
        RECT  4.350 1.440 4.530 3.940 ;
        RECT  4.290 2.770 4.530 3.940 ;
        RECT  2.710 3.700 4.530 3.940 ;
        RECT  2.710 3.700 2.950 4.620 ;
        RECT  1.990 4.380 2.950 4.620 ;
        RECT  4.990 1.670 5.230 2.230 ;
        RECT  4.830 1.990 5.070 3.390 ;
        RECT  4.770 3.200 5.010 4.620 ;
        RECT  4.770 4.380 5.770 4.620 ;
        RECT  5.950 1.460 6.540 1.700 ;
        RECT  5.790 3.010 6.190 3.410 ;
        RECT  5.950 1.460 6.190 4.060 ;
        RECT  5.950 3.820 7.590 4.060 ;
        RECT  5.310 0.980 7.020 1.220 ;
        RECT  5.310 0.980 5.710 1.380 ;
        RECT  6.780 0.980 7.020 2.200 ;
        RECT  6.780 1.960 8.840 2.200 ;
        RECT  5.470 0.980 5.710 2.710 ;
        RECT  8.600 1.960 8.840 3.000 ;
        RECT  8.600 2.760 9.240 3.000 ;
        RECT  5.310 2.470 5.550 3.810 ;
        RECT  5.250 3.580 5.490 4.140 ;
        RECT  9.090 1.590 9.330 2.520 ;
        RECT  9.090 2.280 9.720 2.520 ;
        RECT  6.430 2.440 6.670 3.570 ;
        RECT  6.430 3.330 9.720 3.570 ;
        RECT  9.480 2.280 9.720 3.650 ;
        RECT  9.210 3.250 9.720 3.650 ;
        RECT  7.900 1.100 11.410 1.340 ;
        RECT  7.900 1.020 8.320 1.430 ;
        RECT  11.170 1.100 11.410 1.750 ;
        RECT  11.170 1.510 11.950 1.750 ;
        RECT  11.710 1.510 11.950 2.540 ;
        RECT  10.450 1.650 10.890 2.050 ;
        RECT  10.450 1.650 10.690 3.500 ;
        RECT  10.450 2.930 10.850 3.500 ;
        RECT  10.450 3.260 12.280 3.500 ;
        RECT  8.050 4.230 9.560 4.470 ;
        RECT  10.830 4.230 12.210 4.470 ;
        RECT  7.550 4.350 8.290 4.590 ;
        RECT  9.320 4.380 11.120 4.620 ;
        RECT  11.980 4.380 12.810 4.620 ;
        RECT  13.280 0.980 13.520 1.780 ;
        RECT  12.200 1.540 14.200 1.780 ;
        RECT  13.960 2.360 15.900 2.600 ;
        RECT  10.950 2.310 11.370 2.710 ;
        RECT  11.130 2.310 11.370 3.020 ;
        RECT  12.200 1.540 12.440 3.020 ;
        RECT  11.130 2.780 12.440 3.020 ;
        RECT  13.960 1.540 14.200 3.500 ;
        RECT  12.580 3.260 14.200 3.500 ;
        RECT  9.750 1.640 10.200 2.040 ;
        RECT  9.960 1.640 10.200 4.140 ;
        RECT  9.960 3.740 13.420 3.990 ;
        RECT  13.180 3.740 13.420 4.270 ;
        RECT  9.960 3.740 10.380 4.140 ;
        RECT  17.440 2.010 17.680 4.270 ;
        RECT  13.180 4.030 17.680 4.270 ;
        RECT  19.710 0.980 20.310 1.220 ;
        RECT  19.710 0.980 19.950 2.410 ;
        RECT  19.710 2.170 20.510 2.410 ;
        RECT  20.270 2.170 20.510 3.410 ;
        RECT  20.270 3.170 20.830 3.410 ;
        RECT  20.770 1.590 22.280 1.830 ;
        RECT  20.770 1.590 21.010 2.920 ;
        RECT  22.040 1.590 22.280 4.130 ;
        RECT  21.730 3.890 22.280 4.130 ;
    END
END sdbfb4

MACRO sdbfb2
    CLASS CORE ;
    FOREIGN sdbfb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.406  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.750 2.020 13.380 2.760 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.456  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.760 2.020 19.000 2.960 ;
        RECT  18.540 2.020 19.000 2.530 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.900 1.960 4.140 2.530 ;
        RECT  3.420 2.580 3.920 3.020 ;
        RECT  3.660 2.290 3.920 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.313  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.150 3.550 15.820 3.790 ;
        RECT  15.580 2.530 15.820 3.790 ;
        RECT  15.420 1.880 15.660 2.770 ;
        RECT  14.620 1.880 15.660 2.120 ;
        RECT  14.620 1.460 15.070 2.120 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.275  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.540 2.020 17.300 2.460 ;
        RECT  16.540 1.510 16.780 4.060 ;
        RECT  16.230 1.410 16.680 1.650 ;
        RECT  16.460 1.510 16.780 1.710 ;
        RECT  16.230 0.980 16.470 1.650 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.010 0.640 2.830 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.370 2.180 3.020 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.760 8.380 3.000 ;
        RECT  7.340 2.580 7.950 3.000 ;
        RECT  7.340 2.580 7.940 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.600 5.600 ;
        RECT  18.310 4.400 18.710 5.600 ;
        RECT  17.100 2.980 17.340 5.600 ;
        RECT  15.740 4.520 16.140 5.600 ;
        RECT  14.380 4.710 14.780 5.600 ;
        RECT  13.180 4.710 13.580 5.600 ;
        RECT  11.350 4.710 11.750 5.600 ;
        RECT  8.680 4.710 9.080 5.600 ;
        RECT  6.420 4.710 6.820 5.600 ;
        RECT  3.190 4.180 3.590 5.600 ;
        RECT  0.720 3.550 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.600 0.740 ;
        RECT  18.460 0.000 18.860 0.890 ;
        RECT  16.890 0.000 17.290 1.290 ;
        RECT  15.410 0.000 15.810 1.620 ;
        RECT  13.900 0.000 14.300 1.260 ;
        RECT  11.880 0.000 12.280 1.260 ;
        RECT  7.420 0.000 7.660 1.720 ;
        RECT  3.320 0.000 3.560 1.200 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.430 1.180 1.670 ;
        RECT  0.900 1.430 1.180 2.420 ;
        RECT  1.050 2.530 1.450 2.930 ;
        RECT  1.050 2.180 1.290 3.310 ;
        RECT  0.230 3.070 1.290 3.310 ;
        RECT  0.230 3.070 0.470 4.620 ;
        RECT  1.510 1.700 2.590 1.940 ;
        RECT  2.350 1.920 3.390 2.130 ;
        RECT  2.420 1.920 3.390 2.160 ;
        RECT  2.420 1.920 2.660 3.460 ;
        RECT  1.540 3.260 2.570 3.500 ;
        RECT  1.540 3.260 1.780 4.000 ;
        RECT  2.040 1.010 3.080 1.250 ;
        RECT  2.840 1.010 3.080 1.680 ;
        RECT  4.520 1.050 4.760 1.600 ;
        RECT  2.840 1.440 4.750 1.680 ;
        RECT  4.520 1.050 4.620 3.010 ;
        RECT  4.380 1.440 4.530 3.940 ;
        RECT  4.290 2.770 4.530 3.940 ;
        RECT  2.710 3.700 4.530 3.940 ;
        RECT  2.710 3.700 2.950 4.620 ;
        RECT  1.990 4.380 2.950 4.620 ;
        RECT  4.990 1.670 5.230 2.230 ;
        RECT  4.860 1.990 5.100 3.390 ;
        RECT  4.770 3.200 5.010 4.620 ;
        RECT  4.770 4.380 5.770 4.620 ;
        RECT  5.980 1.460 6.540 1.700 ;
        RECT  5.820 3.010 6.220 3.410 ;
        RECT  5.980 1.460 6.220 4.060 ;
        RECT  5.980 3.820 7.590 4.060 ;
        RECT  5.310 0.980 7.020 1.220 ;
        RECT  5.310 0.980 5.710 1.430 ;
        RECT  6.780 0.980 7.020 2.200 ;
        RECT  6.780 1.960 8.620 2.200 ;
        RECT  8.380 2.200 8.860 2.440 ;
        RECT  8.620 2.200 8.860 2.930 ;
        RECT  5.470 0.980 5.710 2.710 ;
        RECT  8.620 2.690 9.240 2.930 ;
        RECT  5.340 2.470 5.580 3.810 ;
        RECT  5.250 3.580 5.490 4.140 ;
        RECT  9.010 1.510 9.410 1.910 ;
        RECT  9.160 1.510 9.410 2.450 ;
        RECT  9.160 2.210 9.720 2.450 ;
        RECT  6.460 2.440 6.700 3.570 ;
        RECT  9.280 3.250 9.720 3.650 ;
        RECT  6.460 3.330 9.720 3.570 ;
        RECT  9.480 2.210 9.720 3.650 ;
        RECT  9.260 3.330 9.720 3.650 ;
        RECT  7.900 0.980 11.410 1.220 ;
        RECT  7.900 0.980 8.230 1.430 ;
        RECT  11.170 0.980 11.410 1.990 ;
        RECT  11.170 1.750 11.850 1.990 ;
        RECT  11.610 1.750 11.850 2.540 ;
        RECT  11.610 2.130 12.030 2.540 ;
        RECT  10.440 1.570 10.890 1.970 ;
        RECT  10.440 2.930 10.850 3.310 ;
        RECT  10.440 1.570 10.680 3.310 ;
        RECT  10.610 3.260 12.280 3.500 ;
        RECT  8.050 4.230 9.560 4.470 ;
        RECT  10.830 4.230 12.210 4.470 ;
        RECT  7.550 4.350 8.290 4.590 ;
        RECT  9.320 4.380 11.120 4.620 ;
        RECT  11.980 4.380 12.810 4.620 ;
        RECT  13.280 0.980 13.520 1.780 ;
        RECT  12.270 1.540 14.200 1.780 ;
        RECT  13.960 2.360 15.180 2.600 ;
        RECT  10.950 2.270 11.370 2.670 ;
        RECT  11.130 2.270 11.370 3.020 ;
        RECT  12.200 2.710 12.510 2.950 ;
        RECT  12.270 1.540 12.510 2.950 ;
        RECT  11.130 2.780 12.430 3.020 ;
        RECT  13.960 1.540 14.200 3.450 ;
        RECT  12.580 3.210 14.200 3.450 ;
        RECT  9.750 1.570 10.200 1.970 ;
        RECT  15.900 1.890 16.300 2.290 ;
        RECT  9.960 1.570 10.200 4.140 ;
        RECT  9.950 3.740 12.690 3.990 ;
        RECT  9.950 3.740 10.380 4.140 ;
        RECT  12.450 3.900 13.290 4.140 ;
        RECT  13.050 3.900 13.290 4.470 ;
        RECT  14.830 4.030 16.300 4.270 ;
        RECT  16.060 1.890 16.300 4.270 ;
        RECT  13.050 4.230 15.070 4.470 ;
        RECT  17.530 0.980 18.090 1.220 ;
        RECT  17.530 0.980 17.770 1.760 ;
        RECT  17.540 1.520 17.780 2.440 ;
        RECT  17.620 2.240 17.860 2.920 ;
        RECT  17.820 2.680 18.060 3.490 ;
        RECT  19.050 1.280 19.480 1.700 ;
        RECT  18.030 1.460 19.480 1.700 ;
        RECT  18.030 1.460 18.270 2.020 ;
        RECT  19.240 1.280 19.480 4.210 ;
        RECT  19.040 3.810 19.480 4.210 ;
    END
END sdbfb2

MACRO sdbfb1
    CLASS CORE ;
    FOREIGN sdbfb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.406  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.080 2.580 13.940 3.020 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.456  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.980 2.230 18.420 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.910 2.580 4.440 3.020 ;
        RECT  4.200 2.190 4.440 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.133  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.990 3.570 15.620 3.970 ;
        RECT  15.170 2.870 15.620 3.970 ;
        RECT  15.100 1.580 15.340 3.140 ;
        RECT  14.110 1.580 15.340 1.820 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.181  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.300 1.460 16.740 1.900 ;
        RECT  16.380 1.460 16.620 3.970 ;
        RECT  15.730 1.560 16.740 1.800 ;
        RECT  15.730 1.240 15.970 1.800 ;
        END
    END QN
    PIN SC
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.490 0.750 2.890 ;
        RECT  0.120 2.020 0.580 2.890 ;
        END
    END SC
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.200 2.020 2.740 2.460 ;
        END
    END SD
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.900 2.680 8.710 3.080 ;
        RECT  7.900 2.580 8.380 3.080 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.040 5.600 ;
        RECT  17.580 3.760 17.980 5.600 ;
        RECT  15.590 4.710 16.010 5.600 ;
        RECT  13.870 4.710 14.270 5.600 ;
        RECT  11.680 4.710 12.080 5.600 ;
        RECT  9.010 4.710 9.410 5.600 ;
        RECT  6.750 4.710 7.150 5.600 ;
        RECT  3.170 4.400 3.590 5.600 ;
        RECT  0.720 3.720 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.040 0.740 ;
        RECT  18.260 0.000 18.660 0.960 ;
        RECT  17.490 0.000 17.890 0.960 ;
        RECT  14.880 0.000 15.280 1.280 ;
        RECT  12.290 0.000 12.530 1.600 ;
        RECT  7.740 0.000 7.980 1.720 ;
        RECT  3.410 0.000 3.810 1.430 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.310 1.270 1.550 ;
        RECT  1.030 2.090 1.480 2.490 ;
        RECT  1.030 1.310 1.270 3.370 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.510 1.230 1.960 1.630 ;
        RECT  2.980 2.150 3.560 2.390 ;
        RECT  1.720 1.230 1.960 2.970 ;
        RECT  2.980 2.150 3.220 2.970 ;
        RECT  1.530 2.730 3.220 2.970 ;
        RECT  1.530 2.730 1.770 3.460 ;
        RECT  4.610 1.020 5.010 1.420 ;
        RECT  2.290 1.220 2.530 1.780 ;
        RECT  2.290 1.540 3.180 1.780 ;
        RECT  4.610 1.020 4.920 1.910 ;
        RECT  2.960 1.670 4.920 1.910 ;
        RECT  4.680 1.020 4.920 3.550 ;
        RECT  2.150 3.310 4.920 3.550 ;
        RECT  5.160 1.670 5.400 4.620 ;
        RECT  5.160 4.380 6.200 4.620 ;
        RECT  6.210 1.460 6.820 1.700 ;
        RECT  6.210 1.460 6.450 4.060 ;
        RECT  6.210 3.820 7.920 4.060 ;
        RECT  5.560 0.980 7.300 1.220 ;
        RECT  5.560 0.980 5.960 1.420 ;
        RECT  7.060 0.980 7.300 2.200 ;
        RECT  7.060 1.960 8.880 2.200 ;
        RECT  8.640 2.200 9.190 2.440 ;
        RECT  8.950 2.200 9.190 3.000 ;
        RECT  8.950 2.760 9.570 3.000 ;
        RECT  5.640 0.980 5.880 4.130 ;
        RECT  9.340 1.580 9.740 1.990 ;
        RECT  9.490 1.580 9.740 2.520 ;
        RECT  9.490 2.280 10.050 2.520 ;
        RECT  6.710 2.500 6.950 3.570 ;
        RECT  6.710 3.330 10.050 3.570 ;
        RECT  9.810 2.280 10.050 3.650 ;
        RECT  9.590 3.250 10.050 3.650 ;
        RECT  8.230 1.020 11.740 1.260 ;
        RECT  8.230 1.020 8.640 1.430 ;
        RECT  11.500 1.020 11.740 2.050 ;
        RECT  11.500 1.810 12.160 2.050 ;
        RECT  11.920 1.810 12.160 2.540 ;
        RECT  11.920 2.140 12.360 2.540 ;
        RECT  10.770 1.650 11.220 2.050 ;
        RECT  10.770 1.650 11.010 3.500 ;
        RECT  10.770 2.930 11.180 3.500 ;
        RECT  10.770 3.260 12.610 3.500 ;
        RECT  8.380 4.230 9.890 4.470 ;
        RECT  11.160 4.230 12.540 4.470 ;
        RECT  7.870 4.350 8.620 4.590 ;
        RECT  9.650 4.380 11.450 4.620 ;
        RECT  12.310 4.380 13.140 4.620 ;
        RECT  13.410 1.570 13.810 2.080 ;
        RECT  12.600 1.840 13.810 2.080 ;
        RECT  13.570 1.570 13.810 2.340 ;
        RECT  13.570 2.100 14.530 2.340 ;
        RECT  14.290 2.100 14.530 3.500 ;
        RECT  11.280 2.290 11.680 2.690 ;
        RECT  11.420 2.290 11.680 3.020 ;
        RECT  14.290 2.560 14.860 2.960 ;
        RECT  12.600 1.840 12.840 3.020 ;
        RECT  11.420 2.780 12.840 3.020 ;
        RECT  14.290 2.560 14.690 3.500 ;
        RECT  12.910 3.260 14.690 3.500 ;
        RECT  10.080 1.640 10.530 2.040 ;
        RECT  15.660 2.040 16.100 2.440 ;
        RECT  10.290 1.640 10.530 4.140 ;
        RECT  10.280 3.740 13.620 3.990 ;
        RECT  10.280 3.740 10.710 4.140 ;
        RECT  13.380 3.740 13.620 4.470 ;
        RECT  14.510 4.210 16.100 4.450 ;
        RECT  15.860 2.040 16.100 4.450 ;
        RECT  13.380 4.230 14.700 4.470 ;
        RECT  16.410 0.980 17.220 1.220 ;
        RECT  16.980 0.980 17.220 2.320 ;
        RECT  16.860 2.110 17.100 3.410 ;
        RECT  16.860 3.170 17.410 3.410 ;
        RECT  17.460 1.430 18.900 1.670 ;
        RECT  17.460 1.430 17.710 2.620 ;
        RECT  17.410 2.470 17.650 2.930 ;
        RECT  18.660 1.430 18.900 3.890 ;
        RECT  18.310 3.650 18.900 3.890 ;
    END
END sdbfb1

MACRO ora31d4
    CLASS CORE ;
    FOREIGN ora31d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.000 3.180 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.240 2.020 1.620 2.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.080 2.580 2.740 3.020 ;
        RECT  2.080 2.100 2.320 3.020 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.460 3.300 2.300 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.515  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.740 3.310 5.440 3.580 ;
        RECT  3.740 3.140 4.480 3.580 ;
        RECT  4.240 1.770 4.480 3.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.560 4.240 4.800 5.600 ;
        RECT  3.040 4.530 3.440 5.600 ;
        RECT  0.360 3.960 0.600 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  5.010 0.000 5.410 1.060 ;
        RECT  3.230 0.000 3.470 1.160 ;
        RECT  1.700 0.000 1.940 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.240 0.980 2.790 1.220 ;
        RECT  2.240 0.980 2.480 1.780 ;
        RECT  0.890 1.540 2.480 1.780 ;
        RECT  0.120 1.570 0.550 1.970 ;
        RECT  2.990 2.660 4.000 2.900 ;
        RECT  0.120 1.570 0.360 3.660 ;
        RECT  2.990 2.660 3.230 3.660 ;
        RECT  0.120 3.420 3.230 3.660 ;
    END
END ora31d4

MACRO ora31d2
    CLASS CORE ;
    FOREIGN ora31d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.000 3.180 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.240 2.020 1.620 2.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.080 2.580 2.740 3.020 ;
        RECT  2.080 2.100 2.320 3.020 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.910 1.460 3.300 2.380 ;
        RECT  2.860 1.460 3.300 1.900 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.920 3.340 4.420 3.740 ;
        RECT  4.120 1.350 4.420 3.740 ;
        RECT  3.980 2.580 4.420 3.740 ;
        RECT  3.840 1.350 4.420 1.750 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.540 4.470 4.780 5.600 ;
        RECT  2.970 4.530 3.370 5.600 ;
        RECT  0.360 3.960 0.600 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.570 0.000 4.810 1.160 ;
        RECT  3.230 0.000 3.470 1.160 ;
        RECT  1.710 0.000 1.950 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.250 0.980 2.800 1.220 ;
        RECT  2.250 0.980 2.490 1.780 ;
        RECT  0.900 1.540 2.490 1.780 ;
        RECT  0.120 1.570 0.550 1.970 ;
        RECT  0.120 1.570 0.360 3.660 ;
        RECT  3.440 2.780 3.680 3.660 ;
        RECT  0.120 3.420 3.680 3.660 ;
    END
END ora31d2

MACRO ora31d1
    CLASS CORE ;
    FOREIGN ora31d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.000 3.180 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.940 1.620 2.500 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.080 2.580 2.740 3.020 ;
        RECT  2.080 2.100 2.320 3.020 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.910 1.460 3.300 2.380 ;
        RECT  2.860 1.460 3.300 1.900 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.471  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.930 3.340 4.360 3.740 ;
        RECT  4.120 1.430 4.360 3.740 ;
        RECT  3.980 2.580 4.360 3.740 ;
        RECT  3.930 1.430 4.360 1.830 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  2.940 4.530 3.340 5.600 ;
        RECT  0.360 3.960 0.600 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.260 0.000 3.500 1.200 ;
        RECT  1.740 0.000 1.980 1.170 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.280 0.980 2.830 1.220 ;
        RECT  2.280 0.980 2.520 1.650 ;
        RECT  0.890 1.410 2.520 1.650 ;
        RECT  0.120 1.570 0.550 1.970 ;
        RECT  0.120 1.570 0.360 3.660 ;
        RECT  3.440 2.780 3.680 3.660 ;
        RECT  0.120 3.420 3.680 3.660 ;
    END
END ora31d1

MACRO ora311d4
    CLASS CORE ;
    FOREIGN ora311d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.341  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.020 1.060 2.380 ;
        RECT  0.600 2.020 0.840 3.160 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.313  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 2.580 1.570 3.280 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.459  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.960 2.020 2.200 2.920 ;
        RECT  1.740 2.020 2.200 2.380 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.440 1.840 2.740 3.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.080 2.020 3.860 2.460 ;
        END
    END C3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.857  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.250 3.180 6.010 3.420 ;
        RECT  4.230 1.600 6.010 1.840 ;
        RECT  5.100 1.600 5.540 3.420 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.930 4.570 5.330 5.600 ;
        RECT  3.360 4.570 3.760 5.600 ;
        RECT  0.940 4.180 1.180 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.000 0.000 5.400 0.890 ;
        RECT  3.520 0.000 3.920 0.890 ;
        RECT  2.030 0.000 2.430 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.350 1.360 3.080 1.600 ;
        RECT  1.350 1.360 2.200 1.630 ;
        RECT  0.120 1.460 0.550 1.780 ;
        RECT  4.100 2.240 4.340 2.940 ;
        RECT  2.980 2.700 4.340 2.940 ;
        RECT  0.120 1.460 0.360 4.110 ;
        RECT  0.120 3.600 0.570 4.110 ;
        RECT  0.120 3.700 1.660 3.940 ;
        RECT  0.120 3.700 0.580 4.110 ;
        RECT  2.980 2.700 3.220 4.110 ;
        RECT  1.420 3.870 3.220 4.110 ;
    END
END ora311d4

MACRO ora311d2
    CLASS CORE ;
    FOREIGN ora311d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.343  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.020 1.060 2.380 ;
        RECT  0.600 2.020 0.840 3.160 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.331  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.200 2.580 1.600 3.280 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.459  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.960 2.020 2.200 2.920 ;
        RECT  1.740 2.020 2.200 2.380 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.440 1.840 2.740 3.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.080 2.020 3.860 2.460 ;
        END
    END C3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.248  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.310 3.440 4.980 3.680 ;
        RECT  4.740 1.390 4.980 3.680 ;
        RECT  4.520 2.020 4.980 2.460 ;
        RECT  4.370 1.390 4.980 1.630 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  5.100 4.270 5.340 5.600 ;
        RECT  3.600 4.310 3.840 5.600 ;
        RECT  0.970 4.000 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  5.050 0.000 5.450 0.890 ;
        RECT  3.560 0.000 3.960 0.890 ;
        RECT  2.030 0.000 2.430 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.350 1.360 3.080 1.600 ;
        RECT  1.350 1.360 2.200 1.630 ;
        RECT  0.120 1.460 0.550 1.780 ;
        RECT  2.980 2.700 4.460 2.940 ;
        RECT  0.120 1.460 0.360 3.810 ;
        RECT  0.120 3.520 1.730 3.760 ;
        RECT  0.120 3.410 0.570 3.810 ;
        RECT  1.490 3.520 1.730 4.110 ;
        RECT  2.980 2.700 3.220 4.110 ;
        RECT  1.490 3.870 3.220 4.110 ;
    END
END ora311d2

MACRO ora311d1
    CLASS CORE ;
    FOREIGN ora311d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.341  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.020 1.060 2.460 ;
        RECT  0.600 2.020 0.840 3.160 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.333  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.730 1.620 3.580 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.960 2.020 2.200 2.920 ;
        RECT  1.740 2.020 2.200 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.440 1.840 2.740 3.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.080 1.920 3.860 2.160 ;
        RECT  3.420 1.460 3.860 2.160 ;
        END
    END C3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 1.310 4.920 3.650 ;
        RECT  4.220 1.310 4.920 1.630 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.770 3.970 4.010 5.600 ;
        RECT  1.010 4.330 1.250 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.450 0.000 3.850 1.110 ;
        RECT  2.000 0.000 2.400 1.100 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.350 1.360 3.080 1.600 ;
        RECT  1.350 1.360 2.200 1.630 ;
        RECT  0.120 1.460 0.550 1.780 ;
        RECT  2.980 2.580 4.300 2.820 ;
        RECT  0.120 1.460 0.360 4.090 ;
        RECT  0.120 3.410 0.570 4.090 ;
        RECT  2.980 2.580 3.220 4.090 ;
        RECT  0.120 3.850 3.220 4.090 ;
    END
END ora311d1

MACRO ora21d4
    CLASS CORE ;
    FOREIGN ora21d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.060 3.290 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.491  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.460 3.000 2.180 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.508  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.460 3.300 1.900 ;
        RECT  1.990 2.190 3.100 2.430 ;
        RECT  2.860 1.460 3.100 2.430 ;
        RECT  1.990 2.190 2.390 2.650 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.750 3.130 5.450 3.370 ;
        RECT  3.680 1.850 5.450 2.090 ;
        RECT  4.540 1.850 4.980 3.370 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.360 4.570 4.770 5.600 ;
        RECT  2.710 4.570 3.110 5.600 ;
        RECT  0.500 4.010 0.740 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.450 0.000 4.690 1.330 ;
        RECT  3.090 0.000 3.330 1.190 ;
        RECT  1.580 0.000 1.820 1.390 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.850 1.680 2.610 1.920 ;
        RECT  0.140 1.050 0.550 1.450 ;
        RECT  3.270 2.600 3.870 2.840 ;
        RECT  0.140 1.050 0.380 3.770 ;
        RECT  0.140 3.530 1.220 3.770 ;
        RECT  0.980 3.530 1.220 4.060 ;
        RECT  3.270 2.600 3.510 4.060 ;
        RECT  0.980 3.820 3.510 4.060 ;
    END
END ora21d4

MACRO ora21d2
    CLASS CORE ;
    FOREIGN ora21d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.060 3.290 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.491  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.460 3.000 2.180 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.508  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.910 2.260 3.300 2.500 ;
        RECT  2.860 2.020 3.300 2.500 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.224  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.620 1.770 3.860 3.580 ;
        RECT  3.420 3.140 3.660 3.930 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.010 4.570 4.250 5.600 ;
        RECT  2.510 4.580 2.910 5.600 ;
        RECT  0.500 4.010 0.740 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.310 0.000 4.550 1.510 ;
        RECT  2.950 0.000 3.190 1.510 ;
        RECT  1.580 0.000 1.820 1.320 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.850 1.610 2.570 1.850 ;
        RECT  0.140 0.980 0.550 1.380 ;
        RECT  0.140 0.980 0.380 3.770 ;
        RECT  0.140 3.530 1.220 3.770 ;
        RECT  0.980 3.530 1.220 4.060 ;
        RECT  2.930 3.000 3.170 4.060 ;
        RECT  0.980 3.820 3.170 4.060 ;
    END
END ora21d2

MACRO ora21d1
    CLASS CORE ;
    FOREIGN ora21d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.060 3.290 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.440 3.000 2.180 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.506  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.910 2.260 3.300 2.500 ;
        RECT  2.860 2.020 3.300 2.500 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.159  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.580 1.770 3.860 3.580 ;
        RECT  3.420 3.140 3.660 3.930 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  2.520 4.610 2.920 5.600 ;
        RECT  0.480 4.010 0.720 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  2.950 0.000 3.190 1.510 ;
        RECT  1.580 0.000 1.820 1.320 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.850 1.610 2.570 1.850 ;
        RECT  0.140 0.980 0.550 1.380 ;
        RECT  0.140 0.980 0.380 3.770 ;
        RECT  0.140 3.530 1.200 3.770 ;
        RECT  0.960 3.530 1.200 4.060 ;
        RECT  2.940 3.000 3.180 4.060 ;
        RECT  0.960 3.820 3.180 4.060 ;
    END
END ora21d1

MACRO ora211d4
    CLASS CORE ;
    FOREIGN ora211d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.010 1.060 2.670 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.326  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.030 1.620 3.580 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.680 2.020 2.180 2.670 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.660 2.020 3.300 2.810 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.859  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.250 3.130 6.010 3.370 ;
        RECT  4.230 1.600 6.010 1.840 ;
        RECT  5.100 2.580 5.540 3.370 ;
        RECT  5.300 1.600 5.540 3.370 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.930 4.580 5.330 5.600 ;
        RECT  3.290 4.080 3.530 5.600 ;
        RECT  0.740 4.710 1.140 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.000 0.000 5.400 1.030 ;
        RECT  3.620 0.000 4.020 1.070 ;
        RECT  2.280 0.000 2.680 0.930 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.470 1.270 3.250 1.510 ;
        RECT  0.120 1.530 0.550 1.770 ;
        RECT  3.680 2.320 4.380 2.560 ;
        RECT  3.680 2.320 3.920 3.490 ;
        RECT  2.400 3.250 3.920 3.490 ;
        RECT  0.120 1.530 0.360 4.060 ;
        RECT  0.120 3.660 0.550 4.060 ;
        RECT  2.400 3.250 2.640 4.060 ;
        RECT  0.120 3.820 2.640 4.060 ;
    END
END ora211d4

MACRO ora211d2
    CLASS CORE ;
    FOREIGN ora211d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.326  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.840 0.980 2.470 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.326  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.660 1.650 3.120 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.460  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.660 1.970 2.180 2.380 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.780 3.580 ;
        RECT  2.540 2.660 2.780 3.580 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.350  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.510 3.610 4.440 3.850 ;
        RECT  4.200 1.850 4.440 3.850 ;
        RECT  3.980 3.140 4.440 3.850 ;
        RECT  3.810 1.850 4.440 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.360 4.090 4.600 5.600 ;
        RECT  2.740 4.610 3.140 5.600 ;
        RECT  0.820 4.390 1.060 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.470 0.000 4.870 0.890 ;
        RECT  2.810 0.000 3.210 0.920 ;
        RECT  2.030 0.000 2.430 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.350 1.220 2.770 1.460 ;
        RECT  2.530 1.220 2.770 2.420 ;
        RECT  0.120 0.980 0.550 1.310 ;
        RECT  3.020 2.380 3.960 2.620 ;
        RECT  0.120 0.980 0.360 3.650 ;
        RECT  0.120 3.250 0.550 3.650 ;
        RECT  0.120 3.360 1.910 3.650 ;
        RECT  1.510 3.360 1.910 4.060 ;
        RECT  3.020 2.380 3.260 4.060 ;
        RECT  1.510 3.820 3.260 4.060 ;
    END
END ora211d2

MACRO ora211d1
    CLASS CORE ;
    FOREIGN ora211d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.010 1.060 2.470 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.326  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.030 1.620 3.580 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.460  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.240 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.860 3.580 ;
        RECT  2.620 2.410 2.860 3.580 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.250  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.700 4.330 2.020 ;
        RECT  3.900 1.700 4.140 3.980 ;
        RECT  3.420 1.700 4.140 2.460 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.060 4.610 3.460 5.600 ;
        RECT  1.140 4.300 1.380 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.160 0.000 3.560 1.100 ;
        RECT  2.030 0.000 2.430 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.350 1.220 2.890 1.460 ;
        RECT  2.650 1.220 2.890 2.170 ;
        RECT  0.120 0.980 0.550 1.310 ;
        RECT  3.100 3.130 3.660 3.370 ;
        RECT  0.120 0.980 0.360 4.060 ;
        RECT  0.120 3.660 0.550 4.060 ;
        RECT  3.100 3.130 3.340 4.060 ;
        RECT  0.120 3.820 3.340 4.060 ;
    END
END ora211d1

MACRO or04da
    CLASS CORE ;
    FOREIGN or04da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 2.020 0.660 3.010 ;
        RECT  0.140 2.020 0.660 2.520 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.000 1.870 2.650 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.110 2.020 2.660 2.510 ;
        RECT  2.110 1.610 2.350 2.510 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.910 2.390 3.300 3.020 ;
        RECT  2.950 1.930 3.190 3.020 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.490 1.090 8.730 3.110 ;
        RECT  5.160 1.610 8.730 3.110 ;
        RECT  4.560 2.500 8.130 4.330 ;
        RECT  6.880 1.180 7.120 4.330 ;
        RECT  3.990 1.340 5.710 1.620 ;
        RECT  5.470 1.180 5.710 4.330 ;
        RECT  3.830 3.770 8.130 4.010 ;
        RECT  3.990 1.180 4.390 1.620 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  8.490 3.340 8.730 5.600 ;
        RECT  7.170 4.620 7.570 5.600 ;
        RECT  5.870 4.620 6.270 5.600 ;
        RECT  4.570 4.620 4.970 5.600 ;
        RECT  3.130 4.620 3.530 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.570 0.000 7.970 0.980 ;
        RECT  6.060 0.000 6.460 0.980 ;
        RECT  4.650 0.000 5.050 0.980 ;
        RECT  3.250 0.000 3.650 0.980 ;
        RECT  1.570 0.000 1.970 0.890 ;
        RECT  0.230 0.000 0.470 1.630 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 4.140 1.860 4.380 ;
        RECT  0.890 1.130 2.940 1.370 ;
        RECT  2.190 0.990 2.940 1.370 ;
        RECT  0.890 1.130 1.850 1.630 ;
        RECT  2.700 1.220 3.750 1.690 ;
        RECT  3.510 1.220 3.750 2.110 ;
        RECT  3.540 1.860 4.920 2.260 ;
        RECT  3.540 1.860 4.310 3.530 ;
        RECT  0.720 3.290 4.310 3.530 ;
        RECT  0.720 3.290 3.440 3.710 ;
    END
END or04da

MACRO or04d7
    CLASS CORE ;
    FOREIGN or04d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 2.020 0.660 3.010 ;
        RECT  0.120 2.020 0.660 2.520 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.000 1.870 2.650 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.110 2.020 2.660 2.510 ;
        RECT  2.110 1.610 2.350 2.510 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.910 2.390 3.300 3.020 ;
        RECT  2.960 1.630 3.200 3.020 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.876  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.510 2.000 7.530 2.510 ;
        RECT  7.290 1.040 7.530 2.510 ;
        RECT  6.510 1.610 6.750 4.090 ;
        RECT  4.260 1.610 6.750 1.850 ;
        RECT  5.740 1.130 5.980 1.850 ;
        RECT  5.210 1.610 5.450 3.830 ;
        RECT  3.830 3.770 4.800 4.010 ;
        RECT  4.560 1.610 4.800 4.010 ;
        RECT  4.260 1.150 4.500 1.850 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  7.170 4.620 7.570 5.600 ;
        RECT  5.870 4.620 6.270 5.600 ;
        RECT  4.570 4.620 4.970 5.600 ;
        RECT  3.130 4.620 3.530 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.400 0.000 6.800 0.980 ;
        RECT  4.920 0.000 5.320 0.980 ;
        RECT  3.160 0.000 3.560 0.890 ;
        RECT  1.570 0.000 1.970 0.890 ;
        RECT  0.230 0.000 0.470 1.630 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 4.140 1.860 4.380 ;
        RECT  2.190 0.990 2.940 1.230 ;
        RECT  0.890 1.130 2.430 1.370 ;
        RECT  2.700 1.130 3.900 1.370 ;
        RECT  0.890 1.130 1.290 1.630 ;
        RECT  3.190 3.290 3.900 3.530 ;
        RECT  3.660 1.130 3.900 3.530 ;
        RECT  0.720 3.470 3.440 3.710 ;
    END
END or04d7

MACRO or04d4
    CLASS CORE ;
    FOREIGN or04d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.340  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.600 0.890 2.840 ;
        RECT  0.120 2.020 0.500 2.840 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.340  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.180 1.840 1.420 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.830 2.020 2.070 2.920 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.386  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.450 1.840 2.690 3.580 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.670 3.130 5.370 3.370 ;
        RECT  3.600 1.850 5.370 2.090 ;
        RECT  4.540 1.850 4.980 3.370 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.310 4.710 4.710 5.600 ;
        RECT  2.930 4.710 3.330 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.310 0.000 4.710 0.890 ;
        RECT  2.930 0.000 3.330 0.890 ;
        RECT  1.330 0.000 1.730 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 1.330 3.330 1.570 ;
        RECT  3.090 2.380 3.700 2.620 ;
        RECT  3.090 1.330 3.330 4.060 ;
        RECT  0.320 3.820 3.330 4.060 ;
    END
END or04d4

MACRO or04d2
    CLASS CORE ;
    FOREIGN or04d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.340  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.600 0.890 2.840 ;
        RECT  0.120 2.020 0.500 2.840 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.340  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.180 1.840 1.420 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.830 2.020 2.070 2.920 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.386  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.450 1.840 2.690 3.580 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.248  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.660 3.130 4.420 3.370 ;
        RECT  3.980 1.850 4.420 3.370 ;
        RECT  3.610 1.850 4.420 2.090 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.310 4.710 4.710 5.600 ;
        RECT  2.730 4.710 3.130 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.310 0.000 4.710 0.890 ;
        RECT  2.930 0.000 3.330 0.890 ;
        RECT  1.370 0.000 1.770 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.760 1.330 3.330 1.570 ;
        RECT  3.090 2.380 3.700 2.620 ;
        RECT  3.090 1.330 3.330 4.060 ;
        RECT  0.320 3.820 3.330 4.060 ;
    END
END or04d2

MACRO or04d1
    CLASS CORE ;
    FOREIGN or04d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.340  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.600 0.890 2.840 ;
        RECT  0.120 2.020 0.500 2.840 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.340  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.180 1.840 1.420 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.830 2.020 2.070 2.920 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.386  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.450 1.840 2.690 3.580 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.240  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.650 1.460 4.020 3.520 ;
        RECT  3.780 1.140 4.020 3.520 ;
        RECT  3.420 1.460 4.020 1.900 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  2.660 4.710 3.060 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  2.930 0.000 3.330 0.890 ;
        RECT  1.370 0.000 1.770 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.760 1.330 3.180 1.570 ;
        RECT  2.940 1.330 3.180 2.490 ;
        RECT  3.170 2.250 3.410 4.060 ;
        RECT  0.320 3.820 3.410 4.060 ;
    END
END or04d1

MACRO or04d0
    CLASS CORE ;
    FOREIGN or04d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.340  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.660 0.890 2.900 ;
        RECT  0.120 2.020 0.500 2.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.340  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.180 1.840 1.420 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.830 2.020 2.070 2.980 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.386  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.450 1.840 2.690 3.580 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.725  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.460 3.200 3.860 3.520 ;
        RECT  3.620 1.290 3.860 3.520 ;
        RECT  3.420 1.290 3.860 1.900 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  2.540 4.710 2.940 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  2.930 0.000 3.330 0.890 ;
        RECT  1.370 0.000 1.770 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.760 1.330 3.180 1.570 ;
        RECT  2.940 1.330 3.180 2.490 ;
        RECT  2.980 2.250 3.220 4.060 ;
        RECT  0.320 3.820 3.220 4.060 ;
    END
END or04d0

MACRO or03da
    CLASS CORE ;
    FOREIGN or03da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.790 0.800 2.190 ;
        RECT  0.120 1.790 0.500 2.460 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 3.140 1.620 3.580 ;
        RECT  1.160 1.790 1.400 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.700 1.930 2.190 2.460 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.034  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.730 1.230 8.160 1.680 ;
        RECT  7.710 1.260 7.950 4.350 ;
        RECT  2.910 2.510 7.950 2.930 ;
        RECT  4.050 1.260 7.950 2.930 ;
        RECT  6.170 1.180 6.570 2.930 ;
        RECT  5.250 1.260 5.490 4.350 ;
        RECT  4.690 1.180 5.090 2.930 ;
        RECT  3.140 1.260 8.160 1.640 ;
        RECT  3.210 1.180 3.610 1.640 ;
        RECT  2.750 3.940 3.150 4.350 ;
        RECT  2.910 2.510 3.150 4.350 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.150 3.180 7.390 5.600 ;
        RECT  5.810 3.160 6.050 5.600 ;
        RECT  4.610 4.620 5.010 5.600 ;
        RECT  3.390 3.160 3.630 5.600 ;
        RECT  2.190 4.620 2.590 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  6.910 0.000 7.310 1.020 ;
        RECT  5.430 0.000 5.830 1.020 ;
        RECT  3.950 0.000 4.350 0.990 ;
        RECT  2.470 0.000 2.860 0.980 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.260 2.860 1.550 ;
        RECT  2.430 1.260 2.860 2.270 ;
        RECT  2.430 1.880 3.810 2.270 ;
        RECT  2.430 1.260 2.670 3.100 ;
        RECT  1.950 2.700 2.670 3.100 ;
        RECT  0.150 3.640 0.550 4.220 ;
        RECT  1.950 2.700 2.390 4.220 ;
        RECT  0.150 3.820 2.390 4.220 ;
    END
END or03da

MACRO or03d7
    CLASS CORE ;
    FOREIGN or03d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.790 0.740 2.190 ;
        RECT  0.120 1.790 0.500 2.460 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.020 3.140 1.620 3.580 ;
        RECT  1.020 2.190 1.400 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.700 1.970 2.190 2.580 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.948  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.100 2.660 6.590 2.900 ;
        RECT  6.090 1.160 6.590 2.900 ;
        RECT  3.110 1.250 6.590 1.490 ;
        RECT  4.100 2.660 4.340 4.340 ;
        RECT  2.710 3.520 4.340 3.760 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.920 4.080 6.320 5.600 ;
        RECT  4.660 3.260 4.900 5.600 ;
        RECT  3.460 4.620 3.870 5.600 ;
        RECT  2.100 4.560 2.500 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.350 0.000 5.750 0.990 ;
        RECT  3.850 0.000 4.250 0.990 ;
        RECT  2.370 0.000 2.770 1.140 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.510 1.230 1.910 1.730 ;
        RECT  0.150 1.310 2.030 1.550 ;
        RECT  1.510 1.490 2.680 1.730 ;
        RECT  2.440 1.860 5.570 2.260 ;
        RECT  2.440 1.490 2.680 3.100 ;
        RECT  2.150 2.860 2.680 3.100 ;
        RECT  0.150 3.660 0.550 4.060 ;
        RECT  2.150 2.860 2.390 4.060 ;
        RECT  0.150 3.820 2.390 4.060 ;
    END
END or03d7

MACRO or03d4
    CLASS CORE ;
    FOREIGN or03d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.265  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.020 1.060 2.570 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.265  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 2.810 1.620 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.265  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.530 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.800  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.130 3.130 4.890 3.370 ;
        RECT  3.120 1.600 4.890 1.840 ;
        RECT  3.980 1.600 4.420 3.370 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.810 4.710 4.210 5.600 ;
        RECT  2.360 4.710 2.760 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.890 0.000 4.290 0.890 ;
        RECT  2.280 0.000 2.680 0.890 ;
        RECT  0.650 0.000 1.050 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.450 0.550 1.780 ;
        RECT  0.120 1.540 2.710 1.780 ;
        RECT  2.470 1.540 2.710 2.560 ;
        RECT  2.470 2.320 3.260 2.560 ;
        RECT  0.120 1.450 0.360 3.740 ;
        RECT  0.120 3.420 0.550 3.740 ;
    END
END or03d4

MACRO or03d2
    CLASS CORE ;
    FOREIGN or03d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.840 1.060 2.460 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.260 2.600 1.500 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.840 2.180 2.460 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.223  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.190 3.140 3.860 3.580 ;
        RECT  3.620 1.830 3.860 3.580 ;
        RECT  3.250 1.830 3.860 2.070 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.930 4.700 4.330 5.600 ;
        RECT  2.570 4.710 2.970 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.930 0.000 4.330 0.890 ;
        RECT  2.280 0.000 2.680 0.890 ;
        RECT  0.920 0.000 1.320 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.240 0.470 1.560 ;
        RECT  0.120 1.320 2.710 1.560 ;
        RECT  2.470 1.320 2.710 2.620 ;
        RECT  2.470 2.380 3.340 2.620 ;
        RECT  0.120 1.240 0.360 3.530 ;
        RECT  0.120 3.210 0.600 3.530 ;
    END
END or03d2

MACRO or03d1
    CLASS CORE ;
    FOREIGN or03d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.840 1.060 2.460 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.260 2.600 1.500 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.840 2.180 2.460 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 3.310 3.580 ;
        RECT  2.990 1.310 3.230 3.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  2.140 4.710 2.540 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  2.140 0.000 2.540 0.890 ;
        RECT  0.920 0.000 1.320 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.240 0.470 1.560 ;
        RECT  0.120 1.320 2.710 1.560 ;
        RECT  2.470 1.320 2.710 2.900 ;
        RECT  0.120 1.240 0.360 3.530 ;
        RECT  0.120 3.210 0.600 3.530 ;
    END
END or03d1

MACRO or03d0
    CLASS CORE ;
    FOREIGN or03d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.840 1.060 2.460 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.260 2.600 1.500 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.840 2.180 2.460 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.818  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 3.190 3.580 ;
        RECT  2.950 1.310 3.190 3.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  2.110 4.710 2.510 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  2.100 0.000 2.500 0.890 ;
        RECT  0.920 0.000 1.320 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.240 0.470 1.560 ;
        RECT  0.120 1.320 2.710 1.560 ;
        RECT  2.470 1.320 2.710 2.900 ;
        RECT  0.120 1.240 0.360 3.530 ;
        RECT  0.120 3.210 0.600 3.530 ;
    END
END or03d0

MACRO or02da
    CLASS CORE ;
    FOREIGN or02da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.280 1.660 0.680 2.060 ;
        RECT  0.120 2.580 0.520 3.020 ;
        RECT  0.280 1.660 0.520 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 1.620 2.460 ;
        RECT  1.090 1.700 1.540 2.100 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.964  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.430 1.230 7.130 1.730 ;
        RECT  6.730 1.150 7.130 1.730 ;
        RECT  2.020 3.180 6.340 3.680 ;
        RECT  3.430 1.230 6.340 3.680 ;
        RECT  2.410 1.220 5.720 1.640 ;
        RECT  5.320 1.110 5.720 3.680 ;
        RECT  3.840 1.110 4.240 3.680 ;
        RECT  2.570 2.520 6.340 3.680 ;
        RECT  2.410 1.110 2.810 1.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.810 4.200 7.050 5.600 ;
        RECT  5.440 4.140 5.680 5.600 ;
        RECT  4.140 4.010 4.380 5.600 ;
        RECT  2.660 4.010 2.900 5.600 ;
        RECT  1.360 3.270 1.600 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.030 0.000 6.430 0.980 ;
        RECT  4.590 0.000 4.990 0.980 ;
        RECT  3.120 0.000 3.520 0.980 ;
        RECT  1.660 0.000 2.060 0.980 ;
        RECT  0.140 0.000 0.560 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.890 1.130 1.470 1.460 ;
        RECT  0.890 1.220 2.170 1.460 ;
        RECT  1.860 1.220 2.170 2.940 ;
        RECT  1.860 1.880 3.190 2.280 ;
        RECT  1.860 1.880 2.330 2.940 ;
        RECT  0.760 2.700 2.330 2.940 ;
        RECT  0.760 2.700 1.760 3.030 ;
        RECT  0.760 2.700 1.120 4.620 ;
        RECT  0.230 3.260 1.120 4.620 ;
    END
END or02da

MACRO or02d7
    CLASS CORE ;
    FOREIGN or02d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.280 1.660 0.680 2.060 ;
        RECT  0.120 2.580 0.520 3.020 ;
        RECT  0.280 1.660 0.520 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.170 2.020 1.620 2.720 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.968  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.240 1.170 5.800 1.420 ;
        RECT  4.730 2.580 5.540 3.020 ;
        RECT  4.290 1.220 5.470 1.460 ;
        RECT  3.390 2.350 5.210 2.750 ;
        RECT  4.810 1.220 5.210 3.020 ;
        RECT  4.730 2.350 5.130 3.740 ;
        RECT  3.790 1.170 4.440 1.420 ;
        RECT  2.720 1.220 3.940 1.460 ;
        RECT  2.090 3.820 3.790 4.220 ;
        RECT  3.390 2.350 3.790 4.220 ;
        RECT  2.390 1.170 2.860 1.420 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.610 4.270 6.010 5.600 ;
        RECT  4.030 3.080 4.270 5.600 ;
        RECT  2.710 4.620 3.110 5.600 ;
        RECT  1.290 3.480 1.690 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.600 0.000 5.000 0.980 ;
        RECT  3.130 0.000 3.530 0.980 ;
        RECT  1.660 0.000 2.060 0.980 ;
        RECT  0.140 0.000 0.560 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.890 1.130 1.470 1.370 ;
        RECT  1.260 1.220 2.150 1.460 ;
        RECT  1.910 1.700 4.390 2.100 ;
        RECT  1.910 1.220 2.150 3.240 ;
        RECT  0.790 3.000 2.150 3.240 ;
        RECT  0.790 3.000 1.030 4.620 ;
        RECT  0.150 4.380 1.030 4.620 ;
    END
END or02d7

MACRO or02d4
    CLASS CORE ;
    FOREIGN or02d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.120 0.830 2.360 ;
        RECT  0.120 1.460 0.500 2.360 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.170 2.320 1.620 3.020 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.844  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.570 1.850 4.330 2.090 ;
        RECT  2.490 3.130 4.240 3.370 ;
        RECT  3.420 1.850 3.860 3.370 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.150 4.710 3.560 5.600 ;
        RECT  1.750 4.710 2.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.280 0.000 3.680 0.890 ;
        RECT  1.880 0.000 2.280 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 1.540 2.100 1.780 ;
        RECT  1.860 2.380 2.520 2.620 ;
        RECT  1.860 1.540 2.100 3.500 ;
        RECT  0.150 3.260 2.100 3.500 ;
    END
END or02d4

MACRO or02d2
    CLASS CORE ;
    FOREIGN or02d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.810 2.540 ;
        RECT  0.120 1.440 0.500 2.540 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.410 3.580 ;
        RECT  1.170 2.220 1.410 3.580 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.460 2.680 1.900 ;
        RECT  2.300 1.460 2.540 3.700 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.800 4.710 3.200 5.600 ;
        RECT  1.380 4.710 1.780 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.840 0.000 3.210 0.890 ;
        RECT  1.250 0.000 1.650 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 1.720 2.060 1.960 ;
        RECT  1.820 1.720 2.060 4.090 ;
        RECT  0.150 3.850 2.060 4.090 ;
    END
END or02d2

MACRO or02d1
    CLASS CORE ;
    FOREIGN or02d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.810 2.540 ;
        RECT  0.120 1.440 0.500 2.540 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.410 3.580 ;
        RECT  1.170 2.220 1.410 3.580 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.375  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.460 2.680 1.900 ;
        RECT  2.300 1.460 2.570 3.700 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  1.380 4.710 1.780 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  1.290 0.000 1.690 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 1.720 2.060 1.960 ;
        RECT  1.820 1.720 2.060 4.090 ;
        RECT  0.150 3.850 2.060 4.090 ;
    END
END or02d1

MACRO or02d0
    CLASS CORE ;
    FOREIGN or02d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.810 2.540 ;
        RECT  0.120 1.440 0.500 2.540 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.410 3.580 ;
        RECT  1.170 2.220 1.410 3.580 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.718  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.460 2.680 2.090 ;
        RECT  2.300 1.460 2.570 3.700 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  1.380 4.710 1.780 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  1.290 0.000 1.690 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 1.720 2.060 1.960 ;
        RECT  1.820 1.720 2.060 4.090 ;
        RECT  0.150 3.850 2.060 4.090 ;
    END
END or02d0

MACRO oan211d4
    CLASS CORE ;
    FOREIGN oan211d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.460 3.300 2.540 ;
        RECT  2.860 1.460 3.300 1.900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.800 2.480 2.180 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.310 0.500 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.580 3.580 ;
        RECT  1.180 2.170 1.420 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.032  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.810 3.130 6.570 3.370 ;
        RECT  4.810 1.830 6.570 2.070 ;
        RECT  5.660 1.830 6.100 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.490 4.710 5.890 5.600 ;
        RECT  3.990 4.710 4.390 5.600 ;
        RECT  1.380 4.710 1.780 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.550 0.000 5.950 0.890 ;
        RECT  4.150 0.000 4.550 0.890 ;
        RECT  2.810 0.000 3.210 0.890 ;
        RECT  0.770 0.000 1.250 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.690 1.870 1.930 ;
        RECT  1.820 3.260 2.400 3.500 ;
        RECT  1.820 3.260 2.060 4.060 ;
        RECT  0.150 3.820 2.060 4.060 ;
        RECT  2.290 1.610 2.530 2.260 ;
        RECT  2.420 2.040 2.660 3.020 ;
        RECT  3.630 2.520 3.950 3.020 ;
        RECT  2.420 2.780 3.950 3.020 ;
        RECT  2.820 2.780 3.060 3.470 ;
        RECT  3.590 1.730 3.830 2.280 ;
        RECT  3.590 2.040 4.430 2.280 ;
        RECT  4.190 2.360 4.960 2.600 ;
        RECT  4.190 2.040 4.430 3.500 ;
        RECT  3.510 3.260 4.430 3.500 ;
    END
END oan211d4

MACRO oan211d2
    CLASS CORE ;
    FOREIGN oan211d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.460 3.300 2.540 ;
        RECT  2.860 1.460 3.300 1.900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.800 2.480 2.180 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.310 0.500 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.580 3.580 ;
        RECT  1.180 2.170 1.420 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.242  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.810 3.130 5.540 3.450 ;
        RECT  5.300 1.570 5.540 3.450 ;
        RECT  5.100 2.580 5.540 3.450 ;
        RECT  4.870 1.570 5.540 1.810 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.550 4.710 5.950 5.600 ;
        RECT  4.180 4.710 4.580 5.600 ;
        RECT  1.380 4.710 1.780 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.550 0.000 5.950 0.890 ;
        RECT  4.150 0.000 4.550 0.890 ;
        RECT  2.810 0.000 3.210 0.890 ;
        RECT  0.810 0.000 1.210 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.690 1.870 1.930 ;
        RECT  1.820 3.260 2.400 3.500 ;
        RECT  1.820 3.260 2.060 4.060 ;
        RECT  0.150 3.820 2.060 4.060 ;
        RECT  2.290 1.610 2.530 2.260 ;
        RECT  2.420 2.040 2.660 3.020 ;
        RECT  3.630 2.520 3.950 3.020 ;
        RECT  2.420 2.780 3.950 3.020 ;
        RECT  2.820 2.780 3.060 3.470 ;
        RECT  3.590 1.490 3.830 2.060 ;
        RECT  3.590 1.820 4.430 2.060 ;
        RECT  4.190 2.100 4.960 2.340 ;
        RECT  4.190 1.820 4.430 3.500 ;
        RECT  3.510 3.260 4.430 3.500 ;
    END
END oan211d2

MACRO oan211d1
    CLASS CORE ;
    FOREIGN oan211d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.460 3.240 2.520 ;
        RECT  2.860 1.460 3.240 1.900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.800 2.480 2.180 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.310 0.500 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.580 3.580 ;
        RECT  1.180 2.150 1.420 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.132  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.740 3.060 4.140 ;
        RECT  2.820 2.780 3.060 4.140 ;
        RECT  2.420 2.780 3.060 3.020 ;
        RECT  2.420 2.040 2.660 3.020 ;
        RECT  2.290 1.590 2.530 2.260 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  1.460 4.300 1.700 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.890 0.000 3.130 1.220 ;
        RECT  0.890 0.000 1.130 1.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.670 1.870 1.910 ;
        RECT  1.820 3.260 2.400 3.500 ;
        RECT  1.820 3.260 2.060 4.060 ;
        RECT  0.150 3.820 2.060 4.060 ;
    END
END oan211d1

MACRO oaim3m11d4
    CLASS CORE ;
    FOREIGN oaim3m11d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.940 4.150 2.460 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.350 5.540 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.520 1.060 3.020 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 1.900 ;
        RECT  1.270 1.460 1.510 2.330 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.520 2.180 3.020 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.847  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.610 3.130 9.370 3.370 ;
        RECT  7.590 1.600 9.370 1.840 ;
        RECT  8.460 1.600 8.900 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  8.290 4.570 8.690 5.600 ;
        RECT  6.870 4.570 7.270 5.600 ;
        RECT  4.990 4.370 5.230 5.600 ;
        RECT  3.630 3.660 3.870 5.600 ;
        RECT  2.140 4.520 2.540 5.600 ;
        RECT  0.760 4.520 1.160 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.330 0.000 8.730 1.060 ;
        RECT  6.960 0.000 7.360 1.060 ;
        RECT  5.640 0.000 5.880 1.370 ;
        RECT  2.310 0.000 2.550 1.240 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.390 0.550 1.720 ;
        RECT  2.430 1.930 2.840 2.250 ;
        RECT  0.120 1.390 0.360 3.580 ;
        RECT  2.430 1.930 2.670 3.500 ;
        RECT  0.120 3.260 2.670 3.500 ;
        RECT  0.120 3.260 0.470 3.580 ;
        RECT  4.550 0.980 5.180 1.220 ;
        RECT  4.940 0.980 5.180 2.110 ;
        RECT  4.940 1.790 6.020 2.110 ;
        RECT  5.780 1.790 6.020 3.650 ;
        RECT  5.520 3.330 6.020 3.650 ;
        RECT  3.990 1.460 4.630 1.700 ;
        RECT  2.910 3.130 4.630 3.370 ;
        RECT  4.210 3.050 4.630 3.450 ;
        RECT  4.390 1.460 4.630 4.130 ;
        RECT  4.390 3.890 5.790 4.130 ;
        RECT  5.550 3.890 5.790 4.540 ;
        RECT  5.550 4.300 6.100 4.540 ;
        RECT  6.290 1.600 7.180 1.840 ;
        RECT  6.940 2.320 7.740 2.560 ;
        RECT  6.940 1.600 7.180 3.130 ;
        RECT  6.310 2.890 7.180 3.130 ;
        RECT  6.310 2.890 6.550 3.450 ;
    END
END oaim3m11d4

MACRO oaim3m11d2
    CLASS CORE ;
    FOREIGN oaim3m11d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.940 4.150 2.460 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.350 5.540 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.520 1.060 3.020 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 1.900 ;
        RECT  1.270 1.460 1.510 2.330 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.520 2.180 3.020 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.248  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.560 3.140 8.340 3.580 ;
        RECT  8.100 1.850 8.340 3.580 ;
        RECT  7.650 1.850 8.340 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  8.350 4.070 8.590 5.600 ;
        RECT  6.990 4.070 7.230 5.600 ;
        RECT  4.990 4.370 5.230 5.600 ;
        RECT  3.630 3.670 3.870 5.600 ;
        RECT  2.140 4.520 2.540 5.600 ;
        RECT  0.760 4.520 1.160 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  8.410 0.000 8.650 1.610 ;
        RECT  7.050 0.000 7.290 1.580 ;
        RECT  5.660 0.000 5.900 1.330 ;
        RECT  2.310 0.000 2.550 1.240 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.390 0.550 1.720 ;
        RECT  2.430 1.930 2.840 2.250 ;
        RECT  0.120 1.390 0.360 3.580 ;
        RECT  2.430 1.930 2.670 3.500 ;
        RECT  0.120 3.260 2.670 3.500 ;
        RECT  0.120 3.260 0.470 3.580 ;
        RECT  4.550 0.980 5.180 1.220 ;
        RECT  4.940 0.980 5.180 2.110 ;
        RECT  4.940 1.790 6.020 2.110 ;
        RECT  5.780 1.790 6.020 3.650 ;
        RECT  5.560 3.330 6.020 3.650 ;
        RECT  3.990 1.460 4.630 1.700 ;
        RECT  2.910 3.130 4.630 3.370 ;
        RECT  4.210 3.040 4.630 3.450 ;
        RECT  4.390 1.460 4.630 4.130 ;
        RECT  4.390 3.890 5.800 4.130 ;
        RECT  5.560 3.890 5.800 4.510 ;
        RECT  5.560 4.270 6.130 4.510 ;
        RECT  6.290 1.850 7.180 2.090 ;
        RECT  6.940 2.380 7.710 2.620 ;
        RECT  6.940 1.850 7.180 3.610 ;
        RECT  6.260 3.370 7.180 3.610 ;
    END
END oaim3m11d2

MACRO oaim3m11d1
    CLASS CORE ;
    FOREIGN oaim3m11d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.940 4.150 2.460 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.350 5.540 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.520 1.060 3.020 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 1.900 ;
        RECT  1.270 1.460 1.510 2.330 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.520 2.180 3.020 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.401  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 3.130 4.630 3.580 ;
        RECT  4.390 1.460 4.630 3.580 ;
        RECT  3.990 1.460 4.630 1.700 ;
        RECT  2.910 3.130 4.630 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.910 4.710 5.310 5.600 ;
        RECT  3.340 4.710 3.740 5.600 ;
        RECT  2.140 4.710 2.540 5.600 ;
        RECT  0.760 4.710 1.160 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.690 0.000 5.930 1.330 ;
        RECT  2.310 0.000 2.550 1.240 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.390 0.550 1.720 ;
        RECT  2.430 1.930 2.840 2.250 ;
        RECT  0.120 1.390 0.360 3.580 ;
        RECT  2.430 1.930 2.670 3.500 ;
        RECT  0.120 3.260 2.670 3.500 ;
        RECT  0.120 3.260 0.470 3.580 ;
        RECT  4.550 0.980 5.180 1.220 ;
        RECT  4.940 0.980 5.180 2.110 ;
        RECT  4.940 1.790 6.040 2.110 ;
        RECT  5.800 1.790 6.040 3.650 ;
        RECT  5.610 3.330 6.040 3.650 ;
    END
END oaim3m11d1

MACRO oaim31d4
    CLASS CORE ;
    FOREIGN oaim31d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  3.420 2.100 3.730 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.790 0.800 3.110 ;
        RECT  0.120 2.020 0.500 3.110 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 3.140 1.620 3.580 ;
        RECT  1.160 2.100 1.400 3.580 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.380 2.500 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.857  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.930 3.130 7.690 3.370 ;
        RECT  5.910 1.600 7.690 1.840 ;
        RECT  6.780 1.600 7.220 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  6.610 4.570 7.010 5.600 ;
        RECT  5.160 4.710 5.560 5.600 ;
        RECT  4.010 4.470 4.250 5.600 ;
        RECT  2.650 4.230 2.890 5.600 ;
        RECT  1.210 4.300 1.450 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.680 0.000 7.080 0.890 ;
        RECT  5.280 0.000 5.680 0.890 ;
        RECT  2.130 0.000 2.530 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 3.050 1.780 ;
        RECT  2.810 1.540 3.050 3.180 ;
        RECT  1.880 2.940 3.050 3.180 ;
        RECT  0.150 3.600 0.550 4.060 ;
        RECT  1.880 2.940 2.120 4.060 ;
        RECT  0.150 3.820 2.120 4.060 ;
        RECT  3.910 1.570 4.360 1.900 ;
        RECT  4.120 2.400 5.020 2.640 ;
        RECT  4.120 1.570 4.360 3.720 ;
        RECT  3.310 3.480 4.360 3.720 ;
        RECT  4.610 1.600 5.500 1.840 ;
        RECT  5.260 2.320 6.060 2.560 ;
        RECT  5.260 1.600 5.500 3.660 ;
        RECT  4.610 3.420 5.500 3.660 ;
    END
END oaim31d4

MACRO oaim31d2
    CLASS CORE ;
    FOREIGN oaim31d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  3.420 2.100 3.730 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.790 0.800 3.110 ;
        RECT  0.120 2.020 0.500 3.110 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 3.140 1.620 3.580 ;
        RECT  1.160 2.100 1.400 3.580 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.380 2.500 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.251  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.880 3.140 6.660 3.580 ;
        RECT  6.420 1.850 6.660 3.580 ;
        RECT  5.960 1.850 6.660 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.670 4.070 6.910 5.600 ;
        RECT  5.360 4.070 5.600 5.600 ;
        RECT  4.010 4.480 4.250 5.600 ;
        RECT  2.650 4.230 2.890 5.600 ;
        RECT  1.240 4.300 1.480 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.650 0.000 7.050 0.890 ;
        RECT  5.230 0.000 5.630 0.890 ;
        RECT  2.140 0.000 2.540 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 3.050 1.780 ;
        RECT  2.810 1.540 3.050 3.180 ;
        RECT  1.880 2.940 3.050 3.180 ;
        RECT  0.150 3.600 0.550 4.060 ;
        RECT  1.880 2.940 2.120 4.060 ;
        RECT  0.150 3.820 2.120 4.060 ;
        RECT  3.910 1.570 4.360 1.900 ;
        RECT  4.120 2.600 5.020 2.840 ;
        RECT  4.120 1.570 4.360 3.720 ;
        RECT  3.310 3.480 4.360 3.720 ;
        RECT  4.610 1.850 5.500 2.090 ;
        RECT  5.260 2.380 6.030 2.620 ;
        RECT  5.260 1.850 5.500 3.370 ;
        RECT  4.660 3.130 5.500 3.370 ;
        RECT  4.660 3.130 4.900 3.690 ;
    END
END oaim31d2

MACRO oaim31d1
    CLASS CORE ;
    FOREIGN oaim31d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  3.420 2.100 3.730 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.790 0.800 3.110 ;
        RECT  0.120 2.020 0.500 3.110 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 3.140 1.620 3.580 ;
        RECT  1.160 2.100 1.400 3.580 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.380 2.500 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.331  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.310 3.480 4.360 3.720 ;
        RECT  4.120 1.460 4.360 3.720 ;
        RECT  3.930 1.460 4.360 1.900 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.980 4.230 4.220 5.600 ;
        RECT  2.650 4.230 2.890 5.600 ;
        RECT  1.190 4.300 1.430 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  2.120 0.000 2.520 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 3.050 1.780 ;
        RECT  2.810 1.540 3.050 3.180 ;
        RECT  1.880 2.940 3.050 3.180 ;
        RECT  0.150 3.600 0.550 4.060 ;
        RECT  1.880 2.940 2.120 4.060 ;
        RECT  0.150 3.820 2.120 4.060 ;
    END
END oaim31d1

MACRO oaim311d4
    CLASS CORE ;
    FOREIGN oaim311d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.780 1.780 4.020 2.330 ;
        RECT  3.130 1.780 4.020 2.020 ;
        RECT  2.860 1.460 3.360 1.900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.180 2.580 3.860 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.390 0.500 3.020 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.401  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 1.900 ;
        RECT  1.220 1.460 1.460 2.560 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.421  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.550 2.180 3.020 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.782  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.150 3.130 7.850 3.580 ;
        RECT  5.990 1.600 7.690 1.840 ;
        RECT  6.150 3.120 7.160 3.580 ;
        RECT  6.920 1.600 7.160 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  6.850 4.700 7.250 5.600 ;
        RECT  5.380 4.710 5.780 5.600 ;
        RECT  3.520 4.710 3.920 5.600 ;
        RECT  2.060 4.710 2.460 5.600 ;
        RECT  0.750 4.710 1.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  6.680 0.000 7.080 0.890 ;
        RECT  5.220 0.000 5.620 0.890 ;
        RECT  2.100 0.000 2.500 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 0.940 1.780 ;
        RECT  0.700 1.540 0.940 2.240 ;
        RECT  2.420 2.160 2.900 2.480 ;
        RECT  0.740 2.040 0.980 3.500 ;
        RECT  2.420 2.160 2.660 3.500 ;
        RECT  0.150 3.260 2.660 3.500 ;
        RECT  3.890 1.300 4.500 1.540 ;
        RECT  4.260 1.300 4.500 3.580 ;
        RECT  4.260 2.600 5.290 2.840 ;
        RECT  3.070 3.260 4.520 3.500 ;
        RECT  4.260 2.600 4.520 3.580 ;
        RECT  4.200 3.260 4.520 3.580 ;
        RECT  3.070 3.260 3.310 3.970 ;
        RECT  2.750 3.730 3.310 3.970 ;
        RECT  4.740 1.580 4.980 2.190 ;
        RECT  4.740 1.950 5.770 2.190 ;
        RECT  5.530 2.320 6.330 2.560 ;
        RECT  5.530 1.950 5.770 3.370 ;
        RECT  4.850 3.130 5.770 3.370 ;
    END
END oaim311d4

MACRO oaim311d2
    CLASS CORE ;
    FOREIGN oaim311d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.960 1.800 4.200 2.360 ;
        RECT  3.130 1.800 4.200 2.040 ;
        RECT  2.860 1.460 3.360 1.900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.180 2.580 3.860 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.390 0.500 3.020 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.401  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 1.900 ;
        RECT  1.220 1.460 1.460 2.560 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.421  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.550 2.180 3.020 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.140 3.240 7.160 3.480 ;
        RECT  6.780 1.850 7.160 3.480 ;
        RECT  6.140 1.850 7.160 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.730 4.700 7.130 5.600 ;
        RECT  5.350 4.700 5.750 5.600 ;
        RECT  3.590 4.710 3.990 5.600 ;
        RECT  2.060 4.710 2.460 5.600 ;
        RECT  0.750 4.710 1.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.730 0.000 7.130 0.890 ;
        RECT  5.460 0.000 5.860 0.890 ;
        RECT  2.100 0.000 2.500 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 0.940 1.780 ;
        RECT  0.700 1.540 0.940 2.240 ;
        RECT  2.420 2.160 2.900 2.480 ;
        RECT  0.740 2.040 0.980 3.500 ;
        RECT  2.420 2.160 2.660 3.500 ;
        RECT  0.150 3.260 2.660 3.500 ;
        RECT  3.890 1.320 4.680 1.560 ;
        RECT  4.440 1.320 4.680 2.840 ;
        RECT  4.280 2.600 5.420 2.840 ;
        RECT  4.280 2.600 4.520 3.580 ;
        RECT  2.900 3.260 4.520 3.500 ;
        RECT  4.200 3.260 4.520 3.580 ;
        RECT  2.900 3.260 3.140 3.820 ;
        RECT  4.920 1.770 5.160 2.330 ;
        RECT  4.920 2.090 5.900 2.330 ;
        RECT  5.660 2.380 6.290 2.620 ;
        RECT  5.660 2.090 5.900 3.580 ;
        RECT  4.840 3.340 5.900 3.580 ;
    END
END oaim311d2

MACRO oaim311d1
    CLASS CORE ;
    FOREIGN oaim311d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.920 2.580 4.420 3.020 ;
        RECT  3.920 2.150 4.240 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.300 1.460 3.580 2.990 ;
        RECT  2.860 1.460 3.580 1.900 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.390 0.500 3.020 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.401  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 1.900 ;
        RECT  1.220 1.460 1.460 2.560 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.421  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.550 2.180 3.020 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.480 3.260 4.920 3.580 ;
        RECT  4.680 1.220 4.920 3.580 ;
        RECT  4.540 1.220 4.920 1.900 ;
        RECT  3.890 1.220 4.920 1.470 ;
        RECT  2.990 3.260 4.920 3.500 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.840 4.710 4.240 5.600 ;
        RECT  2.140 4.710 2.540 5.600 ;
        RECT  0.750 4.710 1.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  2.180 0.000 2.420 1.540 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 0.940 1.780 ;
        RECT  0.700 1.540 0.940 2.240 ;
        RECT  2.420 2.160 2.900 2.480 ;
        RECT  0.740 2.040 0.980 3.500 ;
        RECT  2.420 2.160 2.660 3.500 ;
        RECT  0.150 3.260 2.660 3.500 ;
    END
END oaim311d1

MACRO oaim2m11d4
    CLASS CORE ;
    FOREIGN oaim2m11d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.380 2.480 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.160 2.600 8.840 3.000 ;
        RECT  8.460 2.020 8.840 3.000 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.620 0.850 2.860 ;
        RECT  0.120 2.020 0.500 2.860 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.385  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 2.020 1.620 2.480 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.220 3.130 7.390 3.450 ;
        RECT  7.050 1.770 7.390 3.450 ;
        RECT  5.620 1.850 7.390 2.090 ;
        RECT  6.970 1.770 7.390 2.090 ;
        RECT  6.220 3.130 6.660 3.580 ;
        RECT  5.690 3.130 7.390 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.690 4.700 8.090 5.600 ;
        RECT  6.300 4.710 6.710 5.600 ;
        RECT  4.950 4.710 5.350 5.600 ;
        RECT  2.910 4.710 3.310 5.600 ;
        RECT  1.490 4.710 1.890 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  8.280 0.000 8.680 0.890 ;
        RECT  6.290 0.000 6.690 0.900 ;
        RECT  4.870 0.000 5.270 0.890 ;
        RECT  1.430 0.000 1.830 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 1.540 2.140 1.780 ;
        RECT  1.900 1.540 2.140 2.890 ;
        RECT  1.780 2.670 2.020 3.440 ;
        RECT  0.890 3.200 2.020 3.440 ;
        RECT  2.380 1.540 3.620 1.780 ;
        RECT  3.730 2.450 4.880 2.690 ;
        RECT  2.380 1.540 2.620 3.520 ;
        RECT  2.270 3.120 2.620 3.520 ;
        RECT  2.270 3.200 3.970 3.440 ;
        RECT  2.270 3.200 2.670 3.520 ;
        RECT  3.730 2.450 3.970 3.520 ;
        RECT  3.570 3.120 3.970 3.520 ;
        RECT  4.270 1.840 5.360 2.080 ;
        RECT  5.120 2.380 5.720 2.620 ;
        RECT  5.120 1.840 5.360 3.370 ;
        RECT  4.270 3.130 5.360 3.370 ;
        RECT  7.630 1.540 8.200 1.780 ;
        RECT  7.630 1.540 7.870 3.610 ;
        RECT  7.630 3.370 8.810 3.610 ;
    END
END oaim2m11d4

MACRO oaim2m11d2
    CLASS CORE ;
    FOREIGN oaim2m11d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.380 2.480 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.600 2.600 8.280 3.000 ;
        RECT  7.900 2.020 8.280 3.000 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.620 0.850 2.860 ;
        RECT  0.120 2.020 0.500 2.860 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.385  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 2.020 1.620 2.480 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.242  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 3.050 6.240 3.580 ;
        RECT  5.980 1.850 6.240 3.580 ;
        RECT  5.630 1.850 6.240 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.080 4.700 7.480 5.600 ;
        RECT  6.310 4.710 6.720 5.600 ;
        RECT  4.960 4.710 5.360 5.600 ;
        RECT  2.910 4.710 3.310 5.600 ;
        RECT  1.490 4.710 1.890 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.850 0.000 8.250 0.890 ;
        RECT  6.320 0.000 6.720 0.890 ;
        RECT  4.900 0.000 5.300 0.890 ;
        RECT  1.430 0.000 1.830 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 1.540 2.140 1.780 ;
        RECT  1.900 1.540 2.140 2.890 ;
        RECT  1.780 2.670 2.020 3.440 ;
        RECT  0.890 3.200 2.020 3.440 ;
        RECT  2.380 1.540 3.620 1.780 ;
        RECT  3.800 2.570 4.850 2.810 ;
        RECT  2.380 1.540 2.620 3.520 ;
        RECT  2.270 3.120 2.620 3.520 ;
        RECT  3.800 2.570 4.040 3.520 ;
        RECT  2.270 3.200 4.040 3.520 ;
        RECT  4.280 1.840 5.330 2.080 ;
        RECT  5.090 2.380 5.730 2.620 ;
        RECT  5.090 1.840 5.330 3.370 ;
        RECT  4.280 3.130 5.330 3.370 ;
        RECT  6.990 1.540 7.640 1.780 ;
        RECT  6.990 1.540 7.230 3.610 ;
        RECT  6.990 3.370 8.250 3.610 ;
    END
END oaim2m11d2

MACRO oaim2m11d1
    CLASS CORE ;
    FOREIGN oaim2m11d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.380 2.480 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 5.170 2.460 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.620 0.850 2.860 ;
        RECT  0.120 2.020 0.500 2.860 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.385  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 2.020 1.620 2.480 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 3.220 3.980 3.460 ;
        RECT  2.380 1.540 3.620 1.780 ;
        RECT  2.270 3.140 2.740 3.580 ;
        RECT  2.380 1.540 2.620 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.280 4.700 4.680 5.600 ;
        RECT  2.710 4.710 3.110 5.600 ;
        RECT  1.490 4.710 1.890 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.890 0.000 5.290 0.890 ;
        RECT  1.430 0.000 1.830 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 1.540 2.140 1.780 ;
        RECT  1.900 1.540 2.140 2.930 ;
        RECT  1.780 2.710 2.020 3.440 ;
        RECT  0.890 3.200 2.020 3.440 ;
        RECT  3.860 1.540 4.660 1.780 ;
        RECT  3.860 1.540 4.100 2.980 ;
        RECT  3.860 2.740 5.340 2.980 ;
        RECT  5.100 2.740 5.340 3.680 ;
    END
END oaim2m11d1

MACRO oaim22d4
    CLASS CORE ;
    FOREIGN oaim22d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.090 2.780 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.700 3.890 2.460 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.720 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 2.200 1.620 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.026  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.430 3.300 7.130 3.540 ;
        RECT  6.220 1.690 6.660 3.540 ;
        RECT  5.790 1.690 6.660 1.930 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.050 4.710 6.450 5.600 ;
        RECT  4.690 4.710 5.090 5.600 ;
        RECT  3.490 4.710 3.890 5.600 ;
        RECT  1.460 4.710 1.860 5.600 ;
        RECT  0.170 4.710 0.570 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.620 0.000 7.020 0.980 ;
        RECT  5.190 0.000 5.590 0.980 ;
        RECT  1.430 0.000 1.670 1.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.470 0.980 1.710 ;
        RECT  0.740 1.470 0.980 1.960 ;
        RECT  0.740 1.720 2.100 1.960 ;
        RECT  1.860 1.720 2.100 3.500 ;
        RECT  0.840 3.260 2.100 3.500 ;
        RECT  2.090 1.000 3.830 1.240 ;
        RECT  2.770 1.530 3.260 1.850 ;
        RECT  4.390 2.520 4.710 2.940 ;
        RECT  3.020 2.700 4.710 2.940 ;
        RECT  3.020 1.530 3.260 3.500 ;
        RECT  2.340 3.260 3.260 3.500 ;
        RECT  2.340 3.260 2.580 3.820 ;
        RECT  4.210 0.980 4.450 2.080 ;
        RECT  4.210 1.840 5.190 2.080 ;
        RECT  4.950 2.470 5.460 2.870 ;
        RECT  4.950 1.840 5.190 3.540 ;
        RECT  4.010 3.300 5.190 3.540 ;
    END
END oaim22d4

MACRO oaim22d2
    CLASS CORE ;
    FOREIGN oaim22d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.090 2.780 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.860 3.880 2.460 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.720 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 2.200 1.620 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.470 3.130 6.600 3.370 ;
        RECT  6.220 1.850 6.600 3.370 ;
        RECT  5.490 1.850 6.600 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  6.170 4.710 6.570 5.600 ;
        RECT  4.810 4.700 5.210 5.600 ;
        RECT  3.490 4.710 3.890 5.600 ;
        RECT  1.460 4.710 1.860 5.600 ;
        RECT  0.170 4.710 0.570 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  6.250 0.000 6.490 1.600 ;
        RECT  4.890 0.000 5.130 1.590 ;
        RECT  1.430 0.000 1.670 1.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.470 0.980 1.710 ;
        RECT  0.740 1.470 0.980 1.960 ;
        RECT  0.740 1.720 2.100 1.960 ;
        RECT  1.860 1.720 2.100 3.500 ;
        RECT  0.840 3.260 2.100 3.500 ;
        RECT  2.090 1.000 3.830 1.240 ;
        RECT  2.770 1.530 3.260 1.850 ;
        RECT  4.350 2.520 4.750 2.940 ;
        RECT  3.020 2.700 4.750 2.940 ;
        RECT  3.020 1.530 3.260 3.500 ;
        RECT  2.340 3.260 3.260 3.500 ;
        RECT  2.340 3.260 2.580 3.820 ;
        RECT  4.130 1.850 5.230 2.090 ;
        RECT  4.990 2.380 5.580 2.620 ;
        RECT  4.990 1.850 5.230 3.420 ;
        RECT  4.040 3.180 5.230 3.420 ;
    END
END oaim22d2

MACRO oaim22d1
    CLASS CORE ;
    FOREIGN oaim22d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.392  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.310 0.500 3.020 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.170 3.150 2.460 ;
        RECT  2.340 2.020 2.740 2.460 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.020 4.360 2.790 ;
        END
    END A2
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.392  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 2.580 1.620 3.020 ;
        RECT  1.160 2.200 1.400 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.759  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.140 3.860 3.580 ;
        RECT  2.500 3.130 3.740 3.370 ;
        RECT  3.500 1.600 3.740 3.580 ;
        RECT  3.150 1.600 3.740 1.840 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.730 4.710 4.110 5.600 ;
        RECT  1.510 4.710 1.910 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  1.750 0.000 1.990 1.240 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.480 2.100 1.720 ;
        RECT  1.860 1.480 2.100 3.500 ;
        RECT  0.870 3.260 2.100 3.500 ;
        RECT  2.410 1.000 4.190 1.240 ;
    END
END oaim22d1

MACRO oaim21d4
    CLASS CORE ;
    FOREIGN oaim21d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.520 2.020 2.760 2.790 ;
        RECT  2.300 2.020 2.760 2.460 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 3.140 0.500 3.580 ;
        RECT  0.120 2.650 0.460 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.392  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 2.020 1.400 2.980 ;
        RECT  0.620 2.020 1.400 2.460 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.860 3.130 6.560 3.370 ;
        RECT  4.790 1.850 6.560 2.090 ;
        RECT  5.640 1.850 6.100 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.490 4.710 5.890 5.600 ;
        RECT  4.120 4.710 4.520 5.600 ;
        RECT  2.790 4.710 3.190 5.600 ;
        RECT  1.160 4.710 1.560 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.480 0.000 5.880 0.890 ;
        RECT  4.060 0.000 4.460 0.890 ;
        RECT  1.380 0.000 1.800 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.880 1.780 ;
        RECT  1.640 2.660 2.160 3.060 ;
        RECT  1.640 1.540 1.880 3.510 ;
        RECT  0.750 3.270 1.880 3.510 ;
        RECT  2.690 1.540 3.240 1.780 ;
        RECT  3.000 2.400 4.050 2.640 ;
        RECT  3.000 1.540 3.240 3.540 ;
        RECT  2.120 3.300 3.240 3.540 ;
        RECT  3.520 1.600 4.530 1.840 ;
        RECT  3.520 1.600 3.760 2.160 ;
        RECT  4.290 2.380 4.890 2.620 ;
        RECT  4.290 1.600 4.530 3.180 ;
        RECT  3.520 2.940 4.530 3.180 ;
        RECT  3.520 2.940 3.760 3.510 ;
    END
END oaim21d4

MACRO oaim21d2
    CLASS CORE ;
    FOREIGN oaim21d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.520 2.020 2.760 2.790 ;
        RECT  2.300 2.020 2.760 2.460 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 3.140 0.500 3.580 ;
        RECT  0.120 2.650 0.460 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.392  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 2.020 1.400 2.980 ;
        RECT  0.620 2.020 1.400 2.460 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.248  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.920 3.130 6.040 3.370 ;
        RECT  5.660 1.850 6.040 3.370 ;
        RECT  4.840 1.850 6.040 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.540 4.710 5.940 5.600 ;
        RECT  4.180 4.710 4.580 5.600 ;
        RECT  2.790 4.710 3.190 5.600 ;
        RECT  1.160 4.710 1.560 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.430 0.000 5.830 0.890 ;
        RECT  4.100 0.000 4.550 0.890 ;
        RECT  1.400 0.000 1.800 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.880 1.780 ;
        RECT  1.640 2.660 2.160 3.060 ;
        RECT  1.640 1.540 1.880 3.510 ;
        RECT  0.750 3.270 1.880 3.510 ;
        RECT  2.690 1.540 3.240 1.780 ;
        RECT  3.000 2.380 4.010 2.620 ;
        RECT  3.000 1.540 3.240 3.540 ;
        RECT  2.120 3.300 3.240 3.540 ;
        RECT  3.480 1.850 4.490 2.090 ;
        RECT  4.250 2.380 4.930 2.620 ;
        RECT  4.250 1.850 4.490 3.180 ;
        RECT  3.580 2.940 4.490 3.180 ;
        RECT  3.580 2.940 3.820 3.510 ;
    END
END oaim21d2

MACRO oaim21d1
    CLASS CORE ;
    FOREIGN oaim21d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.520 2.020 2.760 2.790 ;
        RECT  2.300 2.020 2.760 2.460 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 3.140 0.500 3.580 ;
        RECT  0.120 2.650 0.460 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.392  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 2.020 1.400 2.980 ;
        RECT  0.620 2.020 1.400 2.460 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.024  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.120 3.300 3.240 3.580 ;
        RECT  3.000 1.540 3.240 3.580 ;
        RECT  2.860 3.140 3.240 3.580 ;
        RECT  2.690 1.540 3.240 1.780 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.790 4.710 3.190 5.600 ;
        RECT  1.160 4.710 1.560 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  1.400 0.000 1.800 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.880 1.780 ;
        RECT  1.640 2.660 2.160 3.060 ;
        RECT  1.640 1.540 1.880 3.510 ;
        RECT  0.750 3.270 1.880 3.510 ;
    END
END oaim21d1

MACRO oaim211d4
    CLASS CORE ;
    FOREIGN oaim211d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.460 3.300 2.360 ;
        RECT  2.860 1.460 3.300 1.900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.580 2.900 3.060 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.388  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.940 0.500 2.520 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.080 2.020 1.620 2.500 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.080  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.420 3.410 7.130 3.650 ;
        RECT  5.420 3.140 6.100 3.650 ;
        RECT  5.850 1.450 6.100 3.650 ;
        RECT  5.420 1.450 6.100 1.690 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.050 4.710 6.450 5.600 ;
        RECT  4.650 4.710 5.050 5.600 ;
        RECT  2.780 4.710 3.180 5.600 ;
        RECT  1.560 4.710 1.960 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.700 0.000 7.100 0.990 ;
        RECT  4.710 0.000 5.110 0.980 ;
        RECT  1.560 0.000 1.800 1.150 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.390 2.100 1.630 ;
        RECT  1.860 1.390 2.100 3.050 ;
        RECT  0.810 2.810 2.100 3.050 ;
        RECT  0.810 2.810 1.050 3.640 ;
        RECT  3.290 0.980 3.840 1.220 ;
        RECT  3.600 0.980 3.840 2.840 ;
        RECT  3.520 2.600 4.700 2.840 ;
        RECT  3.520 2.600 3.780 3.670 ;
        RECT  2.100 3.430 3.780 3.670 ;
        RECT  3.540 2.600 3.780 4.070 ;
        RECT  4.080 1.170 4.320 2.140 ;
        RECT  4.080 1.900 5.180 2.140 ;
        RECT  4.940 2.490 5.490 2.890 ;
        RECT  4.940 1.900 5.180 3.370 ;
        RECT  4.080 3.130 5.180 3.370 ;
    END
END oaim211d4

MACRO oaim211d2
    CLASS CORE ;
    FOREIGN oaim211d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.460 3.380 2.360 ;
        RECT  2.860 1.460 3.380 1.900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.580 2.900 3.060 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.388  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.020 0.500 2.720 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.080 2.020 1.620 2.500 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.246  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.760 1.420 6.100 3.020 ;
        RECT  5.570 2.580 5.810 3.650 ;
        RECT  5.420 1.420 6.100 1.660 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  6.120 4.710 6.520 5.600 ;
        RECT  4.720 4.710 5.120 5.600 ;
        RECT  2.780 4.710 3.180 5.600 ;
        RECT  1.540 4.710 1.940 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  6.200 0.000 6.440 1.190 ;
        RECT  4.790 0.000 5.030 1.150 ;
        RECT  1.560 0.000 1.800 1.150 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.390 2.100 1.630 ;
        RECT  1.860 1.390 2.100 3.080 ;
        RECT  0.810 2.840 2.100 3.080 ;
        RECT  0.810 2.840 1.050 3.640 ;
        RECT  3.290 0.980 3.860 1.220 ;
        RECT  3.620 2.600 4.810 2.840 ;
        RECT  3.460 3.270 3.860 3.670 ;
        RECT  3.620 0.980 3.860 3.670 ;
        RECT  2.100 3.430 3.860 3.670 ;
        RECT  4.120 1.330 4.360 2.140 ;
        RECT  4.120 1.900 5.520 2.140 ;
        RECT  5.050 1.900 5.520 2.300 ;
        RECT  5.050 1.900 5.290 3.370 ;
        RECT  4.160 3.130 5.290 3.370 ;
    END
END oaim211d2

MACRO oaim211d1
    CLASS CORE ;
    FOREIGN oaim211d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.460 3.530 2.360 ;
        RECT  2.860 1.460 3.530 1.900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.500 2.900 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.388  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.020 0.500 2.720 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.080 2.020 1.620 2.500 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.824  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.050 4.010 3.580 ;
        RECT  3.770 0.980 4.010 3.580 ;
        RECT  3.290 0.980 4.010 1.220 ;
        RECT  2.100 3.290 4.010 3.530 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  2.810 4.710 3.210 5.600 ;
        RECT  1.530 4.710 1.930 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  1.560 0.000 1.800 1.150 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.390 2.100 1.630 ;
        RECT  1.860 1.390 2.100 3.050 ;
        RECT  0.810 2.810 2.100 3.050 ;
        RECT  0.810 2.810 1.050 3.500 ;
    END
END oaim211d1

MACRO oai322d4
    CLASS CORE ;
    FOREIGN oai322d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.690 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.240 3.140 1.620 3.580 ;
        RECT  1.240 2.520 1.530 3.580 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.890 3.580 ;
        RECT  2.650 2.520 2.890 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.020 2.210 2.630 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.478  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.680 3.860 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.490 2.020 4.980 2.460 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.430 2.020 6.100 2.460 ;
        RECT  5.110 2.770 5.670 3.010 ;
        RECT  5.430 2.020 5.670 3.010 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.533  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.380 2.580 8.620 3.620 ;
        RECT  7.070 2.580 8.620 3.020 ;
        RECT  7.710 1.610 7.950 3.020 ;
        RECT  7.070 2.580 7.310 3.620 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.770 4.710 8.170 5.600 ;
        RECT  6.410 4.710 6.810 5.600 ;
        RECT  4.790 4.620 5.190 5.600 ;
        RECT  1.490 4.710 1.890 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  8.410 0.000 8.810 0.980 ;
        RECT  7.000 0.000 7.380 0.980 ;
        RECT  5.520 0.000 5.760 1.160 ;
        RECT  4.200 0.000 4.440 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.110 1.550 1.350 ;
        RECT  1.310 1.110 1.550 1.780 ;
        RECT  1.310 1.540 2.860 1.780 ;
        RECT  2.620 1.760 3.280 2.000 ;
        RECT  2.140 0.980 3.900 1.220 ;
        RECT  3.580 0.980 3.900 1.860 ;
        RECT  3.580 1.540 5.280 1.780 ;
        RECT  3.580 1.540 3.980 1.860 ;
        RECT  0.740 1.700 1.070 2.100 ;
        RECT  5.910 2.700 6.150 3.600 ;
        RECT  4.880 3.360 6.150 3.600 ;
        RECT  0.740 1.700 1.000 4.060 ;
        RECT  4.880 3.360 5.120 4.060 ;
        RECT  0.150 3.820 5.120 4.060 ;
        RECT  6.180 1.540 6.830 1.780 ;
        RECT  6.590 1.540 6.830 4.080 ;
        RECT  5.530 3.840 6.830 4.080 ;
    END
END oai322d4

MACRO oai322d2
    CLASS CORE ;
    FOREIGN oai322d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.630 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.240 3.140 1.620 3.580 ;
        RECT  1.240 2.520 1.530 3.580 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.890 3.580 ;
        RECT  2.650 2.520 2.890 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.020 2.210 2.630 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.478  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.680 3.860 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.500 2.020 4.980 2.460 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.290 2.200 6.100 2.460 ;
        RECT  5.660 2.020 6.100 2.460 ;
        RECT  5.130 2.690 5.530 3.090 ;
        RECT  5.290 2.200 5.530 3.090 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.742  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.460 1.770 8.170 2.090 ;
        RECT  7.930 1.270 8.170 2.090 ;
        RECT  7.160 2.580 7.780 3.020 ;
        RECT  7.460 1.770 7.780 3.020 ;
        RECT  7.160 2.580 7.400 3.990 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.850 4.710 8.250 5.600 ;
        RECT  6.310 4.710 6.710 5.600 ;
        RECT  4.830 4.620 5.230 5.600 ;
        RECT  1.450 4.710 1.850 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.030 0.000 7.270 1.210 ;
        RECT  5.520 0.000 5.760 1.160 ;
        RECT  4.200 0.000 4.440 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.110 1.550 1.350 ;
        RECT  1.310 1.110 1.550 1.780 ;
        RECT  1.310 1.540 2.860 1.780 ;
        RECT  2.620 1.780 3.280 2.020 ;
        RECT  2.140 0.980 3.900 1.220 ;
        RECT  3.580 0.980 3.900 1.860 ;
        RECT  3.580 1.540 5.280 1.780 ;
        RECT  3.580 1.540 3.980 1.860 ;
        RECT  0.740 1.700 1.070 2.100 ;
        RECT  5.890 2.870 6.130 3.600 ;
        RECT  4.280 3.360 6.130 3.600 ;
        RECT  0.740 1.700 1.000 4.060 ;
        RECT  4.280 3.360 4.520 4.060 ;
        RECT  0.150 3.820 4.520 4.060 ;
        RECT  6.180 1.460 6.610 1.780 ;
        RECT  6.370 2.380 6.920 2.620 ;
        RECT  6.370 1.460 6.610 4.080 ;
        RECT  5.570 3.840 6.610 4.080 ;
    END
END oai322d2

MACRO oai322d1
    CLASS CORE ;
    FOREIGN oai322d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.690 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.240 3.140 1.620 3.580 ;
        RECT  1.240 2.520 1.560 3.580 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.570 2.520 3.300 3.030 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.800 2.020 2.210 2.630 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.478  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.540 3.140 4.420 3.580 ;
        RECT  3.540 2.100 3.780 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.150 2.620 4.980 2.860 ;
        RECT  4.540 2.020 4.980 2.860 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.810 3.100 6.040 3.340 ;
        RECT  5.660 2.580 6.040 3.340 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.150 3.820 3.290 4.060 ;
        RECT  2.300 3.700 2.740 4.140 ;
        RECT  0.740 1.700 1.070 2.100 ;
        RECT  0.740 1.700 1.000 4.060 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.880 4.710 5.280 5.600 ;
        RECT  1.490 4.710 1.880 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.560 0.000 5.800 1.160 ;
        RECT  4.220 0.000 4.460 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.110 1.550 1.350 ;
        RECT  1.310 1.110 1.550 1.780 ;
        RECT  1.310 1.540 2.860 1.780 ;
        RECT  2.620 1.780 3.300 2.020 ;
        RECT  2.150 0.990 3.920 1.230 ;
        RECT  3.600 1.540 5.300 1.780 ;
        RECT  3.600 0.990 3.920 1.860 ;
    END
END oai322d1

MACRO oai321d4
    CLASS CORE ;
    FOREIGN oai321d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.490 2.020 4.980 2.460 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.493  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.580 3.300 3.370 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.385  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.890 3.120 4.420 3.580 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.540 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 3.140 1.620 3.580 ;
        RECT  1.160 2.020 1.400 3.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.438  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 3.020 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.110 3.130 8.810 3.370 ;
        RECT  7.040 1.850 8.810 2.090 ;
        RECT  7.900 1.850 8.340 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.720 4.710 8.130 5.600 ;
        RECT  6.370 4.710 6.770 5.600 ;
        RECT  4.110 4.710 4.510 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.810 0.000 8.050 1.330 ;
        RECT  6.390 0.000 6.630 1.330 ;
        RECT  1.470 0.000 1.870 0.980 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.780 1.070 3.750 1.310 ;
        RECT  2.780 1.070 3.030 1.560 ;
        RECT  0.720 1.320 3.030 1.560 ;
        RECT  4.180 1.020 4.420 1.790 ;
        RECT  3.360 1.550 4.420 1.790 ;
        RECT  3.360 1.550 3.600 2.260 ;
        RECT  2.640 2.020 3.600 2.260 ;
        RECT  4.860 0.980 5.460 1.220 ;
        RECT  5.220 2.450 6.300 2.690 ;
        RECT  5.220 0.980 5.460 4.060 ;
        RECT  2.200 3.820 5.460 4.060 ;
        RECT  5.770 1.600 6.780 1.840 ;
        RECT  5.770 1.600 6.010 2.160 ;
        RECT  6.540 2.380 7.140 2.620 ;
        RECT  5.770 3.050 6.010 3.640 ;
        RECT  6.540 1.600 6.780 3.640 ;
        RECT  5.770 3.400 6.780 3.640 ;
    END
END oai321d4

MACRO oai321d2
    CLASS CORE ;
    FOREIGN oai321d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.490 2.020 4.980 2.460 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.493  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.580 3.300 3.370 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.385  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.890 3.120 4.420 3.580 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.540 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 3.140 1.620 3.580 ;
        RECT  1.160 2.020 1.400 3.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.438  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 3.020 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.242  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.110 3.130 8.280 3.370 ;
        RECT  7.900 1.850 8.280 3.370 ;
        RECT  7.040 1.850 8.280 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.720 4.710 8.130 5.600 ;
        RECT  6.370 4.710 6.770 5.600 ;
        RECT  4.110 4.710 4.510 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.810 0.000 8.050 1.330 ;
        RECT  6.390 0.000 6.630 1.330 ;
        RECT  1.470 0.000 1.870 0.980 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.780 1.070 3.750 1.310 ;
        RECT  2.780 1.070 3.030 1.560 ;
        RECT  0.720 1.320 3.030 1.560 ;
        RECT  4.180 1.020 4.420 1.790 ;
        RECT  3.360 1.550 4.420 1.790 ;
        RECT  3.360 1.550 3.600 2.260 ;
        RECT  2.640 2.020 3.600 2.260 ;
        RECT  4.860 0.980 5.460 1.220 ;
        RECT  5.220 2.440 6.300 2.680 ;
        RECT  5.220 0.980 5.460 4.060 ;
        RECT  2.200 3.820 5.460 4.060 ;
        RECT  5.770 1.600 6.780 1.840 ;
        RECT  5.770 1.600 6.010 2.160 ;
        RECT  6.540 2.380 7.140 2.620 ;
        RECT  5.770 3.050 6.010 3.640 ;
        RECT  6.540 1.600 6.780 3.640 ;
        RECT  5.770 3.400 6.780 3.640 ;
    END
END oai321d2

MACRO oai321d1
    CLASS CORE ;
    FOREIGN oai321d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.490 2.020 4.980 2.460 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.493  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.580 3.300 3.370 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.385  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.890 3.120 4.420 3.580 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.540 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 3.140 1.620 3.580 ;
        RECT  1.160 2.020 1.400 3.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.438  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 3.020 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.602  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.210 3.820 5.460 4.060 ;
        RECT  5.220 0.980 5.460 4.060 ;
        RECT  4.860 0.980 5.460 1.220 ;
        RECT  2.210 3.700 2.740 4.140 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.110 4.560 4.510 5.600 ;
        RECT  0.230 3.870 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  1.470 0.000 1.870 0.980 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.780 1.070 3.750 1.310 ;
        RECT  2.780 1.070 3.030 1.560 ;
        RECT  0.720 1.320 3.030 1.560 ;
        RECT  4.180 1.020 4.420 1.790 ;
        RECT  3.360 1.550 4.420 1.790 ;
        RECT  3.360 1.550 3.600 2.260 ;
        RECT  2.640 2.020 3.600 2.260 ;
    END
END oai321d1

MACRO oai31d4
    CLASS CORE ;
    FOREIGN oai31d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.420 0.460 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.486  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.810 1.620 2.540 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.505  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.170 2.740 3.020 ;
        RECT  1.900 2.170 2.740 2.410 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.495  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.460 3.300 1.900 ;
        RECT  2.980 1.460 3.220 2.490 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.849  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.810 3.130 6.570 3.370 ;
        RECT  4.790 1.800 6.570 2.040 ;
        RECT  5.660 1.800 6.100 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.490 4.710 5.890 5.600 ;
        RECT  4.040 4.710 4.440 5.600 ;
        RECT  2.880 4.710 3.280 5.600 ;
        RECT  0.230 4.020 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.650 0.000 5.890 1.290 ;
        RECT  4.190 0.000 4.430 1.290 ;
        RECT  2.940 0.000 3.340 0.890 ;
        RECT  1.540 0.000 1.940 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.770 1.120 1.330 1.360 ;
        RECT  1.090 1.300 2.100 1.540 ;
        RECT  1.860 1.300 2.100 1.880 ;
        RECT  1.860 1.640 2.560 1.880 ;
        RECT  0.150 1.770 0.470 2.180 ;
        RECT  0.150 1.940 0.940 2.180 ;
        RECT  3.700 2.520 4.020 2.970 ;
        RECT  2.980 2.730 4.020 2.970 ;
        RECT  0.700 1.940 0.940 3.620 ;
        RECT  0.700 3.200 1.470 3.620 ;
        RECT  2.980 2.730 3.220 3.620 ;
        RECT  0.700 3.380 3.220 3.620 ;
        RECT  3.570 1.730 3.810 2.280 ;
        RECT  3.570 2.040 4.500 2.280 ;
        RECT  4.260 2.600 4.940 2.840 ;
        RECT  4.260 2.040 4.500 3.450 ;
        RECT  3.510 3.210 4.500 3.450 ;
        RECT  3.510 3.210 3.750 3.770 ;
    END
END oai31d4

MACRO oai31d2
    CLASS CORE ;
    FOREIGN oai31d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.420 0.500 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.810 1.620 2.530 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.504  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.170 2.740 3.020 ;
        RECT  1.860 2.170 2.740 2.410 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.495  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.460 3.300 1.900 ;
        RECT  2.980 1.460 3.220 2.490 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.251  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.770 3.140 5.540 3.580 ;
        RECT  5.300 1.850 5.540 3.580 ;
        RECT  4.840 1.850 5.540 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.500 4.700 5.900 5.600 ;
        RECT  3.970 4.700 4.370 5.600 ;
        RECT  2.610 4.700 3.010 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.610 0.000 5.850 1.600 ;
        RECT  4.230 0.000 4.470 1.580 ;
        RECT  2.940 0.000 3.340 0.890 ;
        RECT  1.540 0.000 1.940 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.770 1.100 1.330 1.340 ;
        RECT  1.090 1.300 2.100 1.540 ;
        RECT  1.860 1.300 2.100 1.880 ;
        RECT  1.860 1.640 2.560 1.880 ;
        RECT  0.150 1.730 0.470 2.180 ;
        RECT  0.150 1.940 0.980 2.180 ;
        RECT  3.460 2.600 4.050 2.840 ;
        RECT  2.980 2.730 3.700 2.970 ;
        RECT  0.740 1.940 0.980 3.500 ;
        RECT  0.740 3.060 1.140 3.500 ;
        RECT  2.980 2.730 3.220 3.500 ;
        RECT  0.740 3.260 3.220 3.500 ;
        RECT  3.570 1.770 3.810 2.330 ;
        RECT  3.570 2.090 4.530 2.330 ;
        RECT  4.290 2.380 4.940 2.620 ;
        RECT  4.290 2.090 4.530 3.450 ;
        RECT  3.490 3.210 4.530 3.450 ;
    END
END oai31d2

MACRO oai31d1
    CLASS CORE ;
    FOREIGN oai31d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.337  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.500 3.580 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.230 2.220 2.180 2.460 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.230 2.220 1.470 2.900 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.420 2.090 2.660 3.580 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.496  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.040 2.130 3.800 2.370 ;
        RECT  3.420 1.460 3.800 2.370 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.309  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.740 3.140 1.620 3.580 ;
        RECT  0.740 1.630 0.980 3.580 ;
        RECT  0.150 1.630 0.980 1.870 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  2.660 4.090 2.900 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  3.270 0.000 3.670 0.890 ;
        RECT  1.670 0.000 2.070 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 1.150 2.770 1.390 ;
        RECT  2.530 1.150 2.770 1.850 ;
    END
END oai31d1

MACRO oai311d4
    CLASS CORE ;
    FOREIGN oai311d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.920 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 2.000 1.620 2.570 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.940 2.020 2.760 2.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  3.000 2.580 3.860 2.820 ;
        RECT  3.000 1.800 3.240 2.820 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.850 1.460 4.410 2.200 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.824  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.990 3.130 7.690 3.370 ;
        RECT  5.920 1.850 7.690 2.090 ;
        RECT  6.770 1.850 7.230 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  6.600 4.710 7.010 5.600 ;
        RECT  5.250 4.710 5.650 5.600 ;
        RECT  3.600 4.710 4.000 5.600 ;
        RECT  0.810 4.710 1.270 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.690 0.000 6.930 1.330 ;
        RECT  5.270 0.000 5.510 1.330 ;
        RECT  3.870 0.000 4.270 0.980 ;
        RECT  2.080 0.000 2.480 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.390 1.280 3.430 1.520 ;
        RECT  0.150 1.170 0.980 1.410 ;
        RECT  4.100 2.450 5.180 2.690 ;
        RECT  0.740 1.170 0.980 3.410 ;
        RECT  0.150 3.170 2.840 3.410 ;
        RECT  4.100 2.450 4.340 3.500 ;
        RECT  2.600 3.260 4.340 3.500 ;
        RECT  4.650 1.600 5.660 1.840 ;
        RECT  4.650 1.600 4.890 2.160 ;
        RECT  5.420 2.380 6.020 2.620 ;
        RECT  4.650 3.050 4.890 3.640 ;
        RECT  5.420 1.600 5.660 3.640 ;
        RECT  4.650 3.400 5.660 3.640 ;
    END
END oai311d4

MACRO oai311d2
    CLASS CORE ;
    FOREIGN oai311d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.920 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 2.000 1.620 2.570 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.880 2.740 2.460 ;
        RECT  1.940 1.880 2.740 2.120 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  3.000 2.580 3.860 2.820 ;
        RECT  3.000 1.800 3.240 2.820 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.850 1.460 4.420 2.200 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.242  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.000 3.130 7.160 3.370 ;
        RECT  6.780 1.850 7.160 3.370 ;
        RECT  5.930 1.850 7.160 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.620 4.710 7.020 5.600 ;
        RECT  5.260 4.710 5.660 5.600 ;
        RECT  3.600 4.710 4.000 5.600 ;
        RECT  0.810 4.710 1.270 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.700 0.000 6.940 1.590 ;
        RECT  5.280 0.000 5.520 1.360 ;
        RECT  3.870 0.000 4.270 0.980 ;
        RECT  2.080 0.000 2.480 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.390 1.280 3.430 1.520 ;
        RECT  0.150 1.540 0.980 1.780 ;
        RECT  4.100 2.440 5.190 2.680 ;
        RECT  0.740 1.540 0.980 3.410 ;
        RECT  0.150 3.170 2.840 3.410 ;
        RECT  4.100 2.440 4.340 3.500 ;
        RECT  2.600 3.260 4.340 3.500 ;
        RECT  4.660 1.600 5.670 1.840 ;
        RECT  4.660 1.600 4.900 2.160 ;
        RECT  5.430 2.380 6.030 2.620 ;
        RECT  5.430 1.600 5.670 3.370 ;
        RECT  4.580 3.130 5.670 3.370 ;
    END
END oai311d2

MACRO oai311d1
    CLASS CORE ;
    FOREIGN oai311d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.930 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 2.020 1.750 2.570 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.160 2.020 2.740 2.630 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  3.000 2.580 3.860 2.820 ;
        RECT  3.000 1.800 3.240 2.820 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 1.460 4.360 2.330 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.876  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.310 3.580 ;
        RECT  0.150 3.170 2.310 3.410 ;
        RECT  0.740 3.140 2.310 3.410 ;
        RECT  0.740 1.170 0.980 3.410 ;
        RECT  0.150 1.170 0.980 1.410 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.600 4.710 4.000 5.600 ;
        RECT  1.160 4.710 1.560 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.910 0.000 4.310 0.980 ;
        RECT  2.080 0.000 2.480 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.390 1.280 3.430 1.530 ;
    END
END oai311d1

MACRO oai22d4
    CLASS CORE ;
    FOREIGN oai22d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.730 2.330 2.140 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.300 2.700 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.820 2.900 1.440 3.140 ;
        RECT  1.200 2.320 1.440 3.140 ;
        RECT  0.620 3.700 1.060 4.140 ;
        RECT  0.820 2.900 1.060 4.140 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.370 0.500 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.857  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.810 3.130 6.570 3.370 ;
        RECT  4.790 1.600 6.570 1.840 ;
        RECT  5.660 2.580 6.100 3.370 ;
        RECT  5.780 1.600 6.020 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.490 4.710 5.890 5.600 ;
        RECT  4.040 4.710 4.440 5.600 ;
        RECT  2.760 4.710 3.160 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.560 0.000 5.960 0.890 ;
        RECT  4.160 0.000 4.560 0.890 ;
        RECT  0.720 0.000 1.120 1.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.450 1.060 1.860 1.380 ;
        RECT  1.450 1.140 3.190 1.380 ;
        RECT  1.450 1.060 1.690 2.080 ;
        RECT  0.150 1.840 1.690 2.080 ;
        RECT  2.180 1.740 2.620 2.060 ;
        RECT  3.580 2.320 3.820 3.180 ;
        RECT  2.380 2.940 3.820 3.180 ;
        RECT  2.380 1.740 2.620 3.700 ;
        RECT  1.380 3.460 2.620 3.700 ;
        RECT  3.570 1.510 3.810 2.080 ;
        RECT  3.570 1.840 4.380 2.080 ;
        RECT  4.140 2.320 4.940 2.560 ;
        RECT  4.140 1.840 4.380 3.660 ;
        RECT  3.430 3.420 4.380 3.660 ;
    END
END oai22d4

MACRO oai22d2
    CLASS CORE ;
    FOREIGN oai22d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.730 2.330 2.140 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.300 2.700 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.820 2.900 1.440 3.140 ;
        RECT  1.200 2.320 1.440 3.140 ;
        RECT  0.620 3.700 1.060 4.140 ;
        RECT  0.820 2.900 1.060 4.140 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.370 0.500 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.251  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.760 3.140 5.540 3.580 ;
        RECT  5.300 1.850 5.540 3.580 ;
        RECT  4.880 1.850 5.540 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.500 4.700 5.900 5.600 ;
        RECT  4.140 4.700 4.540 5.600 ;
        RECT  2.760 4.710 3.160 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.570 0.000 5.970 0.890 ;
        RECT  4.150 0.000 4.550 0.890 ;
        RECT  0.720 0.000 1.120 1.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.450 1.060 1.860 1.380 ;
        RECT  1.450 1.140 3.190 1.380 ;
        RECT  1.450 1.060 1.690 2.080 ;
        RECT  0.150 1.840 1.690 2.080 ;
        RECT  2.180 1.740 2.620 2.060 ;
        RECT  3.580 2.520 3.820 3.180 ;
        RECT  2.380 2.940 3.820 3.180 ;
        RECT  2.380 1.740 2.620 3.700 ;
        RECT  1.380 3.460 2.620 3.700 ;
        RECT  3.570 1.720 3.810 2.280 ;
        RECT  3.570 2.040 4.380 2.280 ;
        RECT  4.140 2.380 4.910 2.620 ;
        RECT  4.140 2.040 4.380 3.660 ;
        RECT  3.460 3.420 4.380 3.660 ;
    END
END oai22d2

MACRO oai22d1
    CLASS CORE ;
    FOREIGN oai22d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.730 2.330 2.140 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.240 2.700 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.820 2.900 1.440 3.140 ;
        RECT  1.200 2.320 1.440 3.140 ;
        RECT  0.620 3.700 1.060 4.140 ;
        RECT  0.820 2.900 1.060 4.140 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.370 0.500 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.380  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.700 2.740 4.140 ;
        RECT  1.380 3.460 2.620 3.700 ;
        RECT  2.380 1.740 2.620 4.140 ;
        RECT  2.180 1.740 2.620 2.060 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.810 4.710 3.210 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  0.800 0.000 1.040 1.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.450 1.060 1.860 1.380 ;
        RECT  1.450 1.140 3.210 1.380 ;
        RECT  1.450 1.060 1.690 2.080 ;
        RECT  0.150 1.840 1.690 2.080 ;
    END
END oai22d1

MACRO oai222d4
    CLASS CORE ;
    FOREIGN oai222d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.489  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 4.980 2.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.350 2.580 3.820 3.080 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.010 2.000 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.478  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.740 3.360 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.020 1.500 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.498  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.800 0.500 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.523  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.540 3.310 8.240 3.580 ;
        RECT  6.540 3.140 7.280 3.580 ;
        RECT  7.040 1.770 7.280 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.280 4.530 7.680 5.600 ;
        RECT  5.980 4.530 6.380 5.600 ;
        RECT  3.370 4.130 3.610 5.600 ;
        RECT  2.550 4.580 2.950 5.600 ;
        RECT  0.150 4.580 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.810 0.000 8.210 1.060 ;
        RECT  5.930 0.000 6.330 1.060 ;
        RECT  1.460 0.000 1.860 0.980 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 1.340 2.960 1.580 ;
        RECT  3.290 1.140 4.890 1.380 ;
        RECT  1.820 2.050 3.530 2.290 ;
        RECT  3.290 1.140 3.530 2.330 ;
        RECT  3.130 1.930 3.530 2.330 ;
        RECT  3.900 1.770 4.300 2.090 ;
        RECT  4.060 3.330 5.780 3.570 ;
        RECT  5.540 2.330 5.780 3.570 ;
        RECT  4.060 1.770 4.300 3.800 ;
        RECT  2.890 3.560 4.300 3.800 ;
        RECT  2.890 3.560 3.130 4.260 ;
        RECT  1.350 4.020 3.130 4.260 ;
        RECT  5.330 1.850 6.300 2.090 ;
        RECT  6.060 2.660 6.790 2.900 ;
        RECT  6.060 1.850 6.300 4.050 ;
        RECT  5.210 3.810 6.300 4.050 ;
    END
END oai222d4

MACRO oai222d2
    CLASS CORE ;
    FOREIGN oai222d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.489  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 4.980 2.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.350 2.580 3.820 3.080 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.010 2.000 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.478  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.740 3.360 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.020 1.500 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.498  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.800 0.500 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.242  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.670 3.130 7.720 3.370 ;
        RECT  7.340 1.850 7.720 3.370 ;
        RECT  6.600 1.850 7.720 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  7.340 4.070 7.580 5.600 ;
        RECT  6.040 4.070 6.280 5.600 ;
        RECT  3.370 4.130 3.610 5.600 ;
        RECT  2.550 4.580 2.950 5.600 ;
        RECT  0.150 4.580 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  7.370 0.000 7.610 1.590 ;
        RECT  6.010 0.000 6.250 1.580 ;
        RECT  1.460 0.000 1.860 0.980 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 1.330 2.960 1.570 ;
        RECT  2.560 1.330 2.960 1.580 ;
        RECT  3.290 1.140 4.890 1.380 ;
        RECT  3.130 1.960 3.530 2.290 ;
        RECT  3.290 1.140 3.530 2.290 ;
        RECT  1.820 2.050 3.530 2.290 ;
        RECT  3.990 1.770 4.230 2.400 ;
        RECT  4.060 3.330 5.090 3.570 ;
        RECT  4.060 2.180 4.300 3.800 ;
        RECT  2.890 3.560 4.300 3.800 ;
        RECT  2.890 3.560 3.130 4.260 ;
        RECT  1.350 4.020 3.130 4.260 ;
        RECT  4.850 3.330 5.090 4.620 ;
        RECT  4.850 4.380 5.720 4.620 ;
        RECT  5.330 2.380 6.700 2.620 ;
        RECT  5.330 1.760 5.570 3.450 ;
    END
END oai222d2

MACRO oai222d1
    CLASS CORE ;
    FOREIGN oai222d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.489  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 4.920 2.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.350 2.580 3.820 3.080 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.010 2.000 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.478  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.740 3.360 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.020 1.500 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.498  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.800 0.500 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.881  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 3.330 4.810 3.570 ;
        RECT  3.980 3.650 4.420 4.140 ;
        RECT  4.060 3.330 4.420 4.140 ;
        RECT  4.060 1.770 4.300 4.140 ;
        RECT  3.910 1.770 4.300 2.170 ;
        RECT  2.890 3.650 4.420 3.890 ;
        RECT  1.350 4.020 3.130 4.260 ;
        RECT  2.890 3.650 3.130 4.260 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.370 4.130 3.610 5.600 ;
        RECT  2.630 4.580 2.870 5.600 ;
        RECT  0.230 4.580 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  1.460 0.000 1.860 0.980 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 1.330 2.960 1.580 ;
        RECT  3.290 1.140 4.890 1.380 ;
        RECT  3.130 1.940 3.530 2.340 ;
        RECT  3.290 1.140 3.530 2.340 ;
        RECT  1.820 2.050 3.530 2.340 ;
    END
END oai222d1

MACRO oai2222d4
    CLASS CORE ;
    FOREIGN oai2222d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.380  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 3.140 9.980 3.580 ;
        RECT  9.740 2.540 9.980 3.580 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.431  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.700 2.580 11.080 3.580 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.790 2.540 9.350 2.780 ;
        RECT  8.790 2.020 9.030 2.780 ;
        RECT  8.460 2.020 9.030 2.460 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.980 1.730 8.220 2.380 ;
        RECT  7.340 1.730 8.220 1.970 ;
        RECT  7.340 1.460 7.780 1.970 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.412  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.700 1.620 4.140 ;
        RECT  1.300 2.580 1.540 4.140 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.431  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.500 3.390 ;
        END
    END C2
    PIN D1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.429  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.980 2.740 2.540 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.412  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 3.140 3.300 3.580 ;
        RECT  3.020 2.020 3.300 3.580 ;
        END
    END D2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.070  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.880 3.140 5.870 3.450 ;
        RECT  3.880 1.490 5.740 1.730 ;
        RECT  3.880 3.140 4.520 3.580 ;
        RECT  3.880 1.490 4.120 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  10.640 4.620 11.040 5.600 ;
        RECT  8.240 4.620 8.640 5.600 ;
        RECT  6.400 4.710 6.800 5.600 ;
        RECT  4.860 4.620 5.260 5.600 ;
        RECT  3.190 4.620 3.590 5.600 ;
        RECT  0.150 4.620 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  8.810 0.000 9.210 0.980 ;
        RECT  7.420 0.000 7.820 0.890 ;
        RECT  6.130 0.000 6.370 1.100 ;
        RECT  4.860 0.000 5.100 1.130 ;
        RECT  3.560 0.000 3.800 1.130 ;
        RECT  2.230 0.000 2.470 1.130 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.730 1.110 1.130 1.610 ;
        RECT  0.730 1.370 2.800 1.610 ;
        RECT  2.560 1.470 3.140 1.710 ;
        RECT  0.150 1.850 2.060 2.090 ;
        RECT  6.110 2.790 6.670 3.030 ;
        RECT  1.820 1.850 2.060 3.240 ;
        RECT  6.110 2.790 6.350 4.060 ;
        RECT  1.860 3.820 6.350 4.060 ;
        RECT  1.860 3.000 2.100 4.620 ;
        RECT  1.470 4.380 2.100 4.620 ;
        RECT  6.730 1.340 6.970 2.550 ;
        RECT  4.630 2.310 7.150 2.550 ;
        RECT  6.910 2.310 7.150 3.770 ;
        RECT  6.910 3.530 8.110 3.770 ;
        RECT  8.160 1.250 10.470 1.490 ;
        RECT  10.070 1.110 10.470 1.510 ;
        RECT  9.270 1.850 11.050 2.090 ;
        RECT  9.270 1.850 9.670 2.300 ;
        RECT  7.540 2.660 7.780 3.260 ;
        RECT  7.540 3.020 8.780 3.260 ;
        RECT  8.540 3.020 8.780 4.150 ;
        RECT  10.220 1.850 10.460 4.150 ;
        RECT  8.540 3.910 10.460 4.150 ;
    END
END oai2222d4

MACRO oai2222d2
    CLASS CORE ;
    FOREIGN oai2222d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.390  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 2.540 8.940 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.140 2.600 10.520 3.580 ;
        RECT  9.660 2.600 10.520 2.840 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.020 8.070 2.460 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.220 1.840 7.100 2.080 ;
        RECT  6.220 1.460 6.660 2.080 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.200 3.140 1.620 3.580 ;
        RECT  1.280 2.520 1.520 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.330 0.500 3.020 ;
        END
    END C2
    PIN D1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.280 2.020 2.740 2.520 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 3.140 3.300 3.580 ;
        RECT  3.020 2.020 3.300 3.580 ;
        END
    END D2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.325  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 1.310 4.630 1.550 ;
        RECT  3.980 2.580 4.420 3.020 ;
        RECT  3.980 2.580 4.310 3.450 ;
        RECT  3.980 1.310 4.300 3.450 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  9.800 4.710 10.200 5.600 ;
        RECT  7.200 4.710 7.600 5.600 ;
        RECT  4.760 4.710 5.160 5.600 ;
        RECT  3.220 4.710 3.620 5.600 ;
        RECT  0.150 4.710 0.560 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  7.750 0.000 8.150 0.980 ;
        RECT  6.360 0.000 6.760 0.980 ;
        RECT  4.910 0.000 5.310 0.980 ;
        RECT  3.500 0.000 3.900 0.980 ;
        RECT  2.160 0.000 2.560 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 1.240 2.480 1.480 ;
        RECT  2.240 1.300 3.160 1.540 ;
        RECT  0.150 1.850 2.040 2.090 ;
        RECT  1.800 1.850 2.040 2.980 ;
        RECT  1.860 2.740 2.100 4.060 ;
        RECT  5.180 2.520 5.420 4.060 ;
        RECT  1.450 3.820 5.420 4.060 ;
        RECT  4.540 1.840 5.910 2.080 ;
        RECT  5.670 1.230 5.910 3.420 ;
        RECT  5.670 3.180 6.850 3.420 ;
        RECT  9.030 1.110 9.430 1.550 ;
        RECT  7.160 1.310 9.430 1.550 ;
        RECT  8.450 1.850 10.170 2.090 ;
        RECT  6.200 2.520 6.600 2.940 ;
        RECT  6.200 2.700 7.330 2.940 ;
        RECT  7.090 2.700 7.330 3.830 ;
        RECT  9.180 1.850 9.420 3.830 ;
        RECT  7.090 3.590 9.420 3.830 ;
    END
END oai2222d2

MACRO oai2222d1
    CLASS CORE ;
    FOREIGN oai2222d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.390  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 2.540 8.940 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.140 2.600 10.520 3.580 ;
        RECT  9.660 2.600 10.520 2.840 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.020 8.070 2.460 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.220 1.840 7.100 2.080 ;
        RECT  6.220 1.460 6.660 2.080 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.180 2.520 1.520 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.330 0.500 3.020 ;
        END
    END C2
    PIN D1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.250 1.800 2.740 2.460 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 3.140 3.300 3.580 ;
        RECT  3.060 2.020 3.300 3.580 ;
        END
    END D2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 1.310 4.630 1.550 ;
        RECT  3.980 2.580 4.420 3.020 ;
        RECT  3.980 1.310 4.300 3.020 ;
        RECT  3.980 1.310 4.250 3.450 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  9.800 4.710 10.200 5.600 ;
        RECT  7.200 4.710 7.600 5.600 ;
        RECT  4.820 4.710 5.220 5.600 ;
        RECT  3.220 4.670 3.620 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  7.750 0.000 8.150 0.980 ;
        RECT  6.360 0.000 6.760 0.980 ;
        RECT  4.910 0.000 5.310 0.980 ;
        RECT  3.500 0.000 3.900 0.980 ;
        RECT  2.160 0.000 2.560 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 1.240 2.480 1.480 ;
        RECT  2.240 1.300 3.160 1.540 ;
        RECT  0.150 1.850 2.010 2.090 ;
        RECT  1.770 1.850 2.010 2.950 ;
        RECT  1.860 2.710 2.100 4.060 ;
        RECT  5.180 2.520 5.420 4.060 ;
        RECT  1.530 3.820 5.420 4.060 ;
        RECT  4.540 1.840 5.910 2.080 ;
        RECT  5.670 1.230 5.910 3.420 ;
        RECT  5.670 3.180 6.850 3.420 ;
        RECT  9.030 1.110 9.430 1.550 ;
        RECT  7.160 1.310 9.430 1.550 ;
        RECT  8.450 1.850 10.170 2.090 ;
        RECT  6.200 2.520 6.600 2.940 ;
        RECT  6.200 2.700 7.330 2.940 ;
        RECT  7.090 2.700 7.330 3.830 ;
        RECT  9.180 1.850 9.420 3.830 ;
        RECT  7.090 3.590 9.420 3.830 ;
    END
END oai2222d1

MACRO oai221d4
    CLASS CORE ;
    FOREIGN oai221d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.360 4.060 2.690 ;
        RECT  3.420 2.360 3.860 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.495  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.730 2.580 2.120 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.360 2.580 2.830 3.200 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.930 1.400 3.170 ;
        RECT  1.160 1.940 1.400 3.170 ;
        RECT  0.620 2.930 1.060 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.690 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.570  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.920 3.290 7.630 3.530 ;
        RECT  6.780 1.690 7.220 3.530 ;
        RECT  6.460 1.690 7.220 1.930 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  6.690 4.710 7.090 5.600 ;
        RECT  5.330 4.710 5.730 5.600 ;
        RECT  3.310 4.710 3.710 5.600 ;
        RECT  2.610 4.710 3.010 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  7.290 0.000 7.690 0.980 ;
        RECT  5.880 0.000 6.260 0.980 ;
        RECT  0.850 0.000 1.090 1.140 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.450 1.190 3.200 1.430 ;
        RECT  1.450 1.190 1.850 1.700 ;
        RECT  0.150 1.460 1.850 1.700 ;
        RECT  2.150 1.780 3.860 2.020 ;
        RECT  4.200 1.840 4.710 2.160 ;
        RECT  4.470 1.840 4.710 3.210 ;
        RECT  4.100 2.970 4.710 3.210 ;
        RECT  2.360 3.580 4.340 3.820 ;
        RECT  3.920 3.420 4.340 3.820 ;
        RECT  4.100 2.970 4.340 3.820 ;
        RECT  1.380 3.820 2.600 4.060 ;
        RECT  4.980 2.630 6.350 2.870 ;
        RECT  4.980 1.760 5.220 3.690 ;
        RECT  4.620 3.450 5.220 3.690 ;
    END
END oai221d4

MACRO oai221d2
    CLASS CORE ;
    FOREIGN oai221d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.450 4.110 2.690 ;
        RECT  3.420 2.450 3.860 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.495  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.730 2.580 2.120 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.360 2.580 2.830 3.200 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.820 2.020 1.480 2.260 ;
        RECT  0.620 2.930 1.060 3.580 ;
        RECT  0.820 2.020 1.060 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.690 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.876  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.140 3.200 7.160 3.440 ;
        RECT  6.780 1.270 7.160 3.440 ;
        RECT  6.340 1.850 7.160 2.090 ;
        RECT  6.730 1.270 7.160 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.810 4.090 7.050 5.600 ;
        RECT  5.430 4.090 5.670 5.600 ;
        RECT  3.410 4.710 3.810 5.600 ;
        RECT  2.760 4.300 3.000 5.600 ;
        RECT  0.260 4.290 0.500 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  5.590 0.000 5.990 0.990 ;
        RECT  0.850 0.000 1.090 1.140 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.450 1.070 3.150 1.310 ;
        RECT  1.450 1.070 1.850 1.700 ;
        RECT  0.150 1.460 1.850 1.700 ;
        RECT  2.150 1.780 3.860 2.020 ;
        RECT  4.200 1.840 4.710 2.160 ;
        RECT  4.470 1.840 4.710 3.170 ;
        RECT  4.100 2.930 4.710 3.170 ;
        RECT  4.100 2.930 4.340 4.060 ;
        RECT  1.480 3.820 4.340 4.060 ;
        RECT  4.730 1.240 5.300 1.480 ;
        RECT  5.060 2.380 6.170 2.620 ;
        RECT  5.060 1.240 5.300 3.650 ;
        RECT  4.720 3.410 5.300 3.650 ;
    END
END oai221d2

MACRO oai221d1
    CLASS CORE ;
    FOREIGN oai221d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 4.300 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.495  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.140 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 2.580 2.860 3.200 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.940 1.410 3.180 ;
        RECT  1.170 1.940 1.410 3.180 ;
        RECT  0.620 2.940 1.060 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.690 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.976  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.510 3.440 4.920 3.680 ;
        RECT  4.540 1.620 4.920 3.680 ;
        RECT  4.430 1.620 4.920 2.020 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.460 4.710 3.860 5.600 ;
        RECT  2.740 4.710 3.140 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  0.850 0.000 1.090 1.140 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.780 1.000 3.380 1.240 ;
        RECT  1.780 1.000 2.020 1.690 ;
        RECT  0.150 1.450 2.020 1.690 ;
        RECT  2.380 1.710 4.090 1.950 ;
    END
END oai221d1

MACRO oai21d4
    CLASS CORE ;
    FOREIGN oai21d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.750 2.250 2.190 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.060 2.650 1.510 3.020 ;
        RECT  0.620 3.700 1.350 4.140 ;
        RECT  1.060 2.650 1.350 4.140 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.250 0.800 2.570 ;
        RECT  0.120 2.250 0.500 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.857  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.250 3.130 6.010 3.370 ;
        RECT  4.230 1.600 6.010 1.840 ;
        RECT  5.100 1.600 5.540 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.930 4.710 5.330 5.600 ;
        RECT  3.480 4.710 3.880 5.600 ;
        RECT  2.250 4.710 2.650 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.000 0.000 5.400 0.890 ;
        RECT  3.600 0.000 4.000 0.890 ;
        RECT  0.890 0.000 1.130 1.190 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.770 1.860 2.010 ;
        RECT  2.230 1.500 2.680 1.900 ;
        RECT  2.440 2.400 3.340 2.640 ;
        RECT  2.440 1.500 2.680 3.500 ;
        RECT  1.590 3.260 2.680 3.500 ;
        RECT  3.010 1.510 3.250 2.080 ;
        RECT  3.010 1.840 3.820 2.080 ;
        RECT  3.580 2.320 4.380 2.560 ;
        RECT  3.580 1.840 3.820 3.120 ;
        RECT  2.950 2.880 3.820 3.120 ;
        RECT  2.950 2.880 3.190 3.450 ;
    END
END oai21d4

MACRO oai21d2
    CLASS CORE ;
    FOREIGN oai21d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.750 2.250 2.190 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.060 2.650 1.510 3.020 ;
        RECT  0.620 3.700 1.350 4.140 ;
        RECT  1.060 2.650 1.350 4.140 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.250 0.800 2.570 ;
        RECT  0.120 2.250 0.500 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.251  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.200 3.140 4.980 3.580 ;
        RECT  4.740 1.850 4.980 3.580 ;
        RECT  4.280 1.850 4.980 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.940 4.700 5.340 5.600 ;
        RECT  3.580 4.700 3.980 5.600 ;
        RECT  2.250 4.700 2.650 5.600 ;
        RECT  0.150 4.700 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.970 0.000 5.370 0.890 ;
        RECT  3.550 0.000 3.950 0.890 ;
        RECT  0.800 0.000 1.220 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.770 1.860 2.010 ;
        RECT  2.230 1.700 2.680 2.010 ;
        RECT  2.440 2.600 3.340 2.840 ;
        RECT  2.440 1.700 2.680 3.500 ;
        RECT  1.590 3.260 2.680 3.500 ;
        RECT  2.930 1.850 3.820 2.090 ;
        RECT  3.580 2.380 4.350 2.620 ;
        RECT  3.580 1.850 3.820 3.370 ;
        RECT  2.980 3.130 3.820 3.370 ;
        RECT  2.980 3.130 3.220 3.690 ;
    END
END oai21d2

MACRO oai21d1
    CLASS CORE ;
    FOREIGN oai21d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.750 2.250 2.190 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.060 3.740 1.620 4.140 ;
        RECT  1.060 2.650 1.510 3.020 ;
        RECT  1.060 2.650 1.350 4.140 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.250 0.800 2.570 ;
        RECT  0.120 2.250 0.500 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.449  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.260 2.680 4.140 ;
        RECT  2.440 1.500 2.680 4.140 ;
        RECT  2.230 1.500 2.680 1.900 ;
        RECT  1.590 3.260 2.680 3.500 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  2.250 4.700 2.650 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  0.770 0.000 1.240 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.770 1.860 2.010 ;
    END
END oai21d1

MACRO oai211d4
    CLASS CORE ;
    FOREIGN oai211d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.449  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.360 2.520 2.760 2.920 ;
        RECT  2.360 2.020 2.740 2.920 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.200 2.120 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.599  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.820 2.780 1.380 3.020 ;
        RECT  1.140 2.200 1.380 3.020 ;
        RECT  0.620 3.140 1.060 3.580 ;
        RECT  0.820 2.780 1.060 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.581  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.710 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.870 3.130 6.570 3.370 ;
        RECT  4.800 1.850 6.570 2.090 ;
        RECT  5.650 1.850 6.110 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.480 4.570 5.890 5.600 ;
        RECT  4.130 4.570 4.530 5.600 ;
        RECT  2.120 4.710 2.520 5.600 ;
        RECT  0.150 4.620 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.570 0.000 5.810 1.330 ;
        RECT  4.150 0.000 4.390 1.320 ;
        RECT  0.930 0.000 1.330 1.150 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.240 1.070 0.480 1.630 ;
        RECT  0.240 1.390 0.960 1.630 ;
        RECT  0.720 1.600 1.960 1.840 ;
        RECT  2.750 1.310 3.290 1.710 ;
        RECT  3.050 2.400 4.060 2.640 ;
        RECT  3.050 1.310 3.290 3.500 ;
        RECT  1.430 3.260 3.290 3.500 ;
        RECT  1.430 3.260 1.670 4.020 ;
        RECT  3.530 1.600 4.540 1.840 ;
        RECT  3.530 1.600 3.770 2.160 ;
        RECT  4.300 2.380 4.900 2.620 ;
        RECT  4.300 1.600 4.540 3.180 ;
        RECT  3.530 2.940 4.540 3.180 ;
        RECT  3.530 2.940 3.770 3.510 ;
    END
END oai211d4

MACRO oai211d2
    CLASS CORE ;
    FOREIGN oai211d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.441  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.360 2.000 2.810 2.920 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.459  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.200 2.120 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.599  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.820 2.610 1.380 2.850 ;
        RECT  1.140 2.200 1.380 2.850 ;
        RECT  0.620 3.140 1.060 3.580 ;
        RECT  0.820 2.610 1.060 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.581  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.710 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.248  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.970 3.130 6.040 3.370 ;
        RECT  5.660 1.850 6.040 3.370 ;
        RECT  4.890 1.850 6.040 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.590 4.710 5.990 5.600 ;
        RECT  4.230 4.710 4.630 5.600 ;
        RECT  2.080 4.710 2.480 5.600 ;
        RECT  0.150 4.620 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.660 0.000 5.900 1.610 ;
        RECT  4.240 0.000 4.480 1.550 ;
        RECT  0.930 0.000 1.330 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.160 1.150 0.770 1.390 ;
        RECT  0.530 1.150 0.770 1.710 ;
        RECT  0.530 1.470 2.000 1.710 ;
        RECT  1.600 1.470 2.000 1.870 ;
        RECT  2.830 1.360 3.290 1.760 ;
        RECT  3.050 2.380 4.060 2.620 ;
        RECT  1.430 3.260 3.290 3.500 ;
        RECT  3.050 1.360 3.290 3.660 ;
        RECT  2.840 3.260 3.290 3.660 ;
        RECT  1.430 3.260 1.670 4.020 ;
        RECT  3.530 1.850 4.540 2.090 ;
        RECT  4.300 2.380 4.980 2.620 ;
        RECT  4.300 1.850 4.540 3.180 ;
        RECT  3.630 2.940 4.540 3.180 ;
        RECT  3.630 2.940 3.870 3.510 ;
    END
END oai211d2

MACRO oai211d1
    CLASS CORE ;
    FOREIGN oai211d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.444  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 2.020 2.760 3.030 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.230 2.140 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.599  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.820 2.480 1.410 2.720 ;
        RECT  0.620 3.700 1.060 4.140 ;
        RECT  0.820 2.480 1.060 4.140 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.581  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.290 0.500 3.020 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.999  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 3.270 3.240 4.140 ;
        RECT  3.000 1.290 3.240 4.140 ;
        RECT  2.810 1.290 3.240 1.690 ;
        RECT  1.430 3.430 3.240 3.670 ;
        RECT  2.670 3.270 3.240 3.670 ;
        RECT  1.430 3.430 1.670 4.200 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.170 3.990 2.410 5.600 ;
        RECT  0.150 4.620 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  1.010 0.000 1.250 1.380 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.160 1.230 0.770 1.470 ;
        RECT  0.530 1.230 0.770 1.870 ;
        RECT  0.530 1.630 2.000 1.870 ;
    END
END oai211d1

MACRO nr23d4
    CLASS CORE ;
    FOREIGN nr23d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.508  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.180 0.800 2.580 ;
        RECT  0.120 2.180 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.506  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.420 3.010 ;
        RECT  0.620 1.460 1.420 1.900 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.097  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.100 3.700 3.860 4.140 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.863  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.250 3.130 6.010 3.370 ;
        RECT  4.230 1.520 6.010 1.760 ;
        RECT  5.100 2.580 5.540 3.370 ;
        RECT  5.300 1.520 5.540 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.930 4.570 5.330 5.600 ;
        RECT  3.510 4.570 3.910 5.600 ;
        RECT  1.530 3.940 1.770 5.600 ;
        RECT  0.230 3.940 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.000 0.000 5.400 0.890 ;
        RECT  3.600 0.000 4.000 0.890 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.140 1.620 2.910 1.860 ;
        RECT  2.140 1.620 2.380 3.010 ;
        RECT  2.140 2.770 3.180 3.010 ;
        RECT  2.940 2.770 3.180 3.450 ;
        RECT  1.660 1.130 3.990 1.370 ;
        RECT  3.750 1.130 3.990 2.560 ;
        RECT  3.750 2.320 4.380 2.560 ;
        RECT  1.660 1.130 1.900 3.490 ;
        RECT  0.860 3.250 2.560 3.490 ;
    END
END nr23d4

MACRO nr23d2
    CLASS CORE ;
    FOREIGN nr23d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.508  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.330 0.820 2.570 ;
        RECT  0.120 2.330 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.506  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.420 3.010 ;
        RECT  0.620 1.460 1.420 1.900 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  3.420 2.150 3.660 3.020 ;
        RECT  3.000 2.150 3.660 2.390 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.310 2.580 4.980 3.450 ;
        RECT  4.740 1.620 4.980 3.450 ;
        RECT  4.390 1.620 4.980 1.860 ;
        RECT  4.390 1.300 4.630 1.860 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  5.130 4.130 5.370 5.600 ;
        RECT  3.650 4.130 3.890 5.600 ;
        RECT  1.530 3.940 1.770 5.600 ;
        RECT  0.230 3.940 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  5.130 0.000 5.370 1.250 ;
        RECT  3.540 0.000 3.940 0.890 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.140 1.620 2.910 1.860 ;
        RECT  2.140 1.620 2.380 3.010 ;
        RECT  2.140 2.770 3.180 3.010 ;
        RECT  2.940 2.770 3.180 3.450 ;
        RECT  1.660 1.130 4.140 1.370 ;
        RECT  3.900 1.130 4.140 2.340 ;
        RECT  3.900 2.100 4.500 2.340 ;
        RECT  1.660 1.130 1.900 3.490 ;
        RECT  0.860 3.250 2.560 3.490 ;
    END
END nr23d2

MACRO nr23d1
    CLASS CORE ;
    FOREIGN nr23d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.460 0.770 2.860 ;
        RECT  0.120 2.020 0.500 2.860 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.178  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.580 4.360 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.522  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.180 3.580 ;
        RECT  1.740 1.740 2.020 3.580 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.934  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.260 3.250 1.500 ;
        RECT  2.420 3.080 2.970 3.480 ;
        RECT  2.420 1.260 2.740 3.480 ;
        RECT  2.300 1.260 2.740 1.900 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.530 4.510 3.930 5.600 ;
        RECT  0.860 4.510 1.260 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.680 0.000 3.920 1.440 ;
        RECT  2.260 0.000 2.660 0.930 ;
        RECT  0.880 0.000 1.280 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.280 0.470 1.780 ;
        RECT  0.150 1.540 1.250 1.780 ;
        RECT  1.010 2.500 1.500 2.900 ;
        RECT  1.010 1.540 1.250 3.370 ;
        RECT  0.150 3.130 1.250 3.370 ;
        RECT  3.430 1.850 4.060 2.090 ;
        RECT  2.980 2.600 3.670 2.840 ;
        RECT  3.430 1.850 3.670 3.450 ;
    END
END nr23d1

MACRO nr13d4
    CLASS CORE ;
    FOREIGN nr13d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.504  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 3.010 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.180 0.800 2.500 ;
        RECT  0.120 2.180 0.500 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.580 4.980 3.020 ;
        RECT  3.930 2.580 4.980 2.820 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.996  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.690 1.460 6.570 1.700 ;
        RECT  4.860 3.260 6.560 3.500 ;
        RECT  5.660 1.460 6.100 3.500 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.450 4.580 5.850 5.600 ;
        RECT  4.120 4.580 4.520 5.600 ;
        RECT  2.100 4.710 2.500 5.600 ;
        RECT  0.850 4.510 1.090 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.510 0.000 5.750 1.200 ;
        RECT  3.920 0.000 4.320 0.890 ;
        RECT  0.800 0.000 1.200 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.400 1.780 ;
        RECT  1.160 1.540 1.400 2.980 ;
        RECT  0.740 2.740 1.400 2.980 ;
        RECT  0.740 2.740 0.980 3.500 ;
        RECT  0.150 3.260 0.980 3.500 ;
        RECT  2.900 1.620 3.720 1.860 ;
        RECT  2.900 1.620 3.140 3.370 ;
        RECT  2.900 3.130 3.910 3.370 ;
        RECT  2.420 1.000 2.890 1.370 ;
        RECT  2.420 1.130 4.200 1.370 ;
        RECT  3.960 1.130 4.200 2.340 ;
        RECT  3.960 2.100 5.020 2.340 ;
        RECT  1.530 3.250 2.660 3.500 ;
        RECT  2.420 1.000 2.660 4.050 ;
        RECT  2.420 3.810 3.270 4.050 ;
    END
END nr13d4

MACRO nr13d2
    CLASS CORE ;
    FOREIGN nr13d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.505  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 3.010 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.180 0.800 2.500 ;
        RECT  0.120 2.180 0.500 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.580 4.980 3.020 ;
        RECT  4.090 2.580 4.980 2.820 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.232  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.020 3.260 6.040 3.500 ;
        RECT  5.660 1.460 6.040 3.500 ;
        RECT  4.870 1.460 6.040 1.700 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.610 4.710 6.010 5.600 ;
        RECT  4.250 4.710 4.650 5.600 ;
        RECT  2.280 4.710 2.680 5.600 ;
        RECT  1.000 4.510 1.240 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.690 0.000 5.930 1.200 ;
        RECT  4.100 0.000 4.500 0.890 ;
        RECT  0.800 0.000 1.200 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.400 1.780 ;
        RECT  1.160 1.540 1.400 3.500 ;
        RECT  0.150 3.260 1.400 3.500 ;
        RECT  2.900 1.620 3.750 1.860 ;
        RECT  2.900 1.620 3.140 2.880 ;
        RECT  2.900 2.640 3.850 2.880 ;
        RECT  3.610 2.640 3.850 3.450 ;
        RECT  3.610 3.130 4.080 3.450 ;
        RECT  2.420 1.000 2.890 1.370 ;
        RECT  2.420 1.130 4.230 1.370 ;
        RECT  3.990 1.130 4.230 2.230 ;
        RECT  3.990 1.990 5.170 2.230 ;
        RECT  2.420 1.000 2.660 3.490 ;
        RECT  1.670 3.250 3.370 3.490 ;
    END
END nr13d2

MACRO nr13d1
    CLASS CORE ;
    FOREIGN nr13d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.238  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.070 0.800 2.470 ;
        RECT  0.120 2.070 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.598  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.600 2.470 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.599  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 3.200 3.580 ;
        RECT  2.960 2.520 3.200 3.580 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.554  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.440 1.460 3.680 3.450 ;
        RECT  2.860 1.460 3.680 1.900 ;
        RECT  1.910 1.460 3.680 1.700 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  1.190 4.710 1.590 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  2.530 0.000 2.930 0.890 ;
        RECT  1.170 0.000 1.570 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.500 1.780 ;
        RECT  1.260 1.540 1.500 3.500 ;
        RECT  0.150 3.260 1.500 3.500 ;
    END
END nr13d1

MACRO nr04da
    CLASS CORE ;
    FOREIGN nr04da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.471  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.160 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.471  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.790 2.090 1.350 2.490 ;
        RECT  0.620 2.580 1.060 3.020 ;
        RECT  0.790 2.090 1.060 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.570 2.180 3.020 ;
        RECT  1.740 1.990 1.990 3.020 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.500 2.580 3.220 3.020 ;
        RECT  2.500 2.000 2.740 3.020 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.620 1.240 9.370 2.810 ;
        RECT  4.540 2.570 8.680 4.170 ;
        RECT  5.090 1.190 6.720 1.710 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  8.970 3.080 9.370 5.600 ;
        RECT  7.800 4.620 8.200 5.600 ;
        RECT  6.500 4.620 6.900 5.600 ;
        RECT  5.200 4.620 5.600 5.600 ;
        RECT  3.900 4.620 4.300 5.600 ;
        RECT  2.410 4.100 2.810 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.390 0.000 8.790 0.980 ;
        RECT  7.070 0.000 7.470 0.980 ;
        RECT  5.750 0.000 6.150 0.960 ;
        RECT  4.130 0.000 4.530 0.980 ;
        RECT  2.870 0.000 3.270 1.280 ;
        RECT  1.330 0.000 1.730 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.230 1.130 2.500 1.370 ;
        RECT  2.100 1.030 2.500 1.440 ;
        RECT  2.260 1.030 2.500 1.760 ;
        RECT  0.740 1.310 1.470 1.550 ;
        RECT  2.260 1.520 3.410 1.760 ;
        RECT  3.170 1.520 3.410 2.340 ;
        RECT  3.170 1.940 3.700 2.340 ;
        RECT  3.450 1.940 3.700 3.700 ;
        RECT  1.860 3.460 3.700 3.700 ;
        RECT  0.120 3.620 0.550 4.060 ;
        RECT  1.860 3.460 2.100 4.060 ;
        RECT  0.120 3.820 2.100 4.060 ;
        RECT  3.650 1.290 4.310 1.710 ;
        RECT  3.930 1.940 5.390 2.340 ;
        RECT  3.930 1.290 4.310 4.360 ;
        RECT  3.130 3.960 4.310 4.360 ;
    END
END nr04da

MACRO nr04d7
    CLASS CORE ;
    FOREIGN nr04d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.650 2.920 ;
        RECT  0.120 2.020 0.500 2.920 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.150 3.220 1.620 3.580 ;
        RECT  1.150 1.860 1.390 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.180 2.940 ;
        RECT  1.830 1.840 2.070 2.940 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 2.660 3.300 2.940 ;
        RECT  2.510 2.660 3.300 2.900 ;
        RECT  2.510 2.110 2.750 2.900 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.596  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.250 2.600 8.130 2.840 ;
        RECT  7.730 1.420 8.130 2.840 ;
        RECT  5.080 1.480 8.130 1.660 ;
        RECT  6.960 1.420 8.130 1.660 ;
        RECT  7.320 2.600 7.560 4.240 ;
        RECT  7.250 2.600 7.560 3.900 ;
        RECT  5.300 3.660 7.560 3.900 ;
        RECT  6.780 3.140 7.560 3.900 ;
        RECT  6.050 1.480 7.130 1.720 ;
        RECT  4.620 1.420 6.250 1.590 ;
        RECT  4.640 3.840 5.660 4.080 ;
        RECT  4.280 1.350 5.370 1.460 ;
        RECT  4.280 1.220 4.840 1.460 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.850 3.150 8.250 5.600 ;
        RECT  6.680 4.620 7.080 5.600 ;
        RECT  5.380 4.620 5.780 5.600 ;
        RECT  4.070 4.620 4.470 5.600 ;
        RECT  2.340 3.810 2.960 4.050 ;
        RECT  2.340 3.810 2.580 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.850 0.000 8.250 1.160 ;
        RECT  6.440 0.000 6.840 1.210 ;
        RECT  4.960 0.000 5.360 1.010 ;
        RECT  2.840 1.110 3.390 1.350 ;
        RECT  3.150 0.000 3.390 1.350 ;
        RECT  1.330 0.000 1.730 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.100 1.030 2.500 1.550 ;
        RECT  0.740 1.310 2.600 1.550 ;
        RECT  2.360 1.310 2.600 1.860 ;
        RECT  2.360 1.620 3.230 1.860 ;
        RECT  2.990 1.620 3.230 2.420 ;
        RECT  2.990 2.180 3.860 2.420 ;
        RECT  3.620 2.180 3.860 3.570 ;
        RECT  1.860 3.330 3.860 3.570 ;
        RECT  0.290 3.170 0.530 4.060 ;
        RECT  1.860 3.330 2.100 4.060 ;
        RECT  0.290 3.820 2.100 4.060 ;
        RECT  3.660 1.380 3.900 1.940 ;
        RECT  3.660 1.700 4.380 1.940 ;
        RECT  4.140 2.120 7.490 2.360 ;
        RECT  4.140 1.700 4.380 4.050 ;
        RECT  3.300 3.810 4.380 4.050 ;
    END
END nr04d7

MACRO nr04d4
    CLASS CORE ;
    FOREIGN nr04d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.330 0.800 2.730 ;
        RECT  0.120 1.460 0.500 2.730 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 3.140 1.620 3.580 ;
        RECT  1.160 2.520 1.400 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.840 2.020 2.080 2.970 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.760 3.580 ;
        RECT  2.520 2.690 2.760 3.580 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.853  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.810 3.130 6.570 3.370 ;
        RECT  4.800 1.600 6.510 1.840 ;
        RECT  5.660 1.600 6.100 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.490 4.710 5.890 5.600 ;
        RECT  4.030 4.710 4.430 5.600 ;
        RECT  2.740 4.710 3.140 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.570 0.000 5.970 0.890 ;
        RECT  4.180 0.000 4.580 0.890 ;
        RECT  2.800 0.000 3.200 0.890 ;
        RECT  1.170 0.000 1.570 0.890 ;
        RECT  0.230 0.000 0.630 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.260 1.540 3.240 1.780 ;
        RECT  1.260 1.540 1.500 2.090 ;
        RECT  0.820 1.850 1.500 2.090 ;
        RECT  3.000 2.400 3.920 2.640 ;
        RECT  3.000 1.540 3.240 4.060 ;
        RECT  0.150 3.820 3.240 4.060 ;
        RECT  3.580 1.510 3.820 2.080 ;
        RECT  3.580 1.840 4.400 2.080 ;
        RECT  4.160 2.320 4.960 2.560 ;
        RECT  4.160 1.840 4.400 3.120 ;
        RECT  3.520 2.880 4.400 3.120 ;
        RECT  3.520 2.880 3.760 3.740 ;
    END
END nr04d4

MACRO nr04d2
    CLASS CORE ;
    FOREIGN nr04d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.330 0.800 2.730 ;
        RECT  0.120 1.460 0.500 2.730 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 3.140 1.620 3.580 ;
        RECT  1.160 2.520 1.400 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.840 2.020 2.080 2.970 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.760 3.580 ;
        RECT  2.520 2.690 2.760 3.580 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.251  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.780 3.140 5.560 3.580 ;
        RECT  5.320 1.850 5.560 3.580 ;
        RECT  4.900 1.850 5.560 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.520 4.700 5.920 5.600 ;
        RECT  4.160 4.700 4.560 5.600 ;
        RECT  2.740 4.710 3.140 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.590 0.000 5.990 0.890 ;
        RECT  4.170 0.000 4.570 0.890 ;
        RECT  2.810 0.000 3.210 0.890 ;
        RECT  1.180 0.000 1.580 0.890 ;
        RECT  0.230 0.000 0.630 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.260 1.540 3.240 1.780 ;
        RECT  1.260 1.540 1.500 2.090 ;
        RECT  0.820 1.850 1.500 2.090 ;
        RECT  3.000 2.600 3.920 2.840 ;
        RECT  3.000 1.540 3.240 4.060 ;
        RECT  0.150 3.820 3.240 4.060 ;
        RECT  3.590 1.720 3.830 2.280 ;
        RECT  3.590 2.040 4.400 2.280 ;
        RECT  4.160 2.380 4.930 2.620 ;
        RECT  4.160 2.040 4.400 3.660 ;
        RECT  3.480 3.420 4.400 3.660 ;
    END
END nr04d2

MACRO nr04d1
    CLASS CORE ;
    FOREIGN nr04d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.760 3.580 ;
        RECT  2.520 2.690 2.760 3.580 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.840 2.020 2.080 2.970 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 3.140 1.620 3.580 ;
        RECT  1.160 2.520 1.400 3.580 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.330 0.800 2.730 ;
        RECT  0.120 1.460 0.500 2.730 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.824  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.150 3.820 3.240 4.060 ;
        RECT  3.000 1.540 3.240 4.060 ;
        RECT  2.860 1.540 3.240 2.460 ;
        RECT  1.260 1.540 3.240 1.780 ;
        RECT  0.820 1.850 1.500 2.090 ;
        RECT  1.260 1.540 1.500 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.740 4.710 3.140 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.810 0.000 3.210 0.890 ;
        RECT  1.180 0.000 1.580 0.890 ;
        RECT  0.230 0.000 0.630 0.890 ;
        END
    END VSS
END nr04d1

MACRO nr04d0
    CLASS CORE ;
    FOREIGN nr04d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.243  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.760 3.580 ;
        RECT  2.520 2.690 2.760 3.580 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.243  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.460 ;
        RECT  1.840 2.020 2.080 2.970 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.243  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 3.140 1.620 3.580 ;
        RECT  1.160 2.570 1.400 3.580 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.243  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.110 0.800 2.510 ;
        RECT  0.120 1.460 0.500 2.510 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.974  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.150 3.820 3.240 4.060 ;
        RECT  3.000 1.540 3.240 4.060 ;
        RECT  2.860 1.540 3.240 2.460 ;
        RECT  1.320 1.540 3.240 1.780 ;
        RECT  0.830 1.600 1.560 1.840 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.740 4.710 3.140 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.810 0.000 3.210 0.890 ;
        RECT  1.180 0.000 1.580 0.890 ;
        RECT  0.230 0.000 0.630 0.890 ;
        END
    END VSS
END nr04d0

MACRO nr03da
    CLASS CORE ;
    FOREIGN nr03da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.610 2.350 1.060 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.467  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.690 1.620 4.140 ;
        RECT  1.350 1.980 1.620 4.140 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.467  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.040 3.080 2.660 3.600 ;
        RECT  2.040 2.260 2.280 3.600 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.954  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.930 2.280 9.400 4.350 ;
        RECT  4.880 2.280 9.400 2.900 ;
        RECT  4.880 1.220 8.620 2.900 ;
        RECT  8.220 1.080 8.620 2.900 ;
        RECT  6.740 1.080 7.140 2.900 ;
        RECT  6.300 1.220 6.800 4.350 ;
        RECT  3.880 2.510 6.800 3.010 ;
        RECT  3.860 1.130 5.660 1.620 ;
        RECT  5.260 1.080 5.660 3.010 ;
        RECT  3.880 2.510 4.380 4.380 ;
        RECT  3.860 1.080 4.180 1.620 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  8.380 3.180 8.700 5.600 ;
        RECT  7.040 3.160 7.440 5.600 ;
        RECT  5.920 4.620 6.320 5.600 ;
        RECT  4.930 3.240 5.170 5.600 ;
        RECT  4.620 3.240 5.170 3.480 ;
        RECT  3.500 4.620 3.900 5.600 ;
        RECT  2.020 4.620 2.420 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.960 0.000 9.360 0.980 ;
        RECT  7.480 0.000 7.880 0.980 ;
        RECT  6.000 0.000 6.400 0.980 ;
        RECT  4.520 0.000 4.920 0.900 ;
        RECT  2.390 0.000 2.630 1.330 ;
        RECT  0.260 1.020 0.820 1.260 ;
        RECT  0.260 0.000 0.500 1.260 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.160 1.010 2.130 1.250 ;
        RECT  1.160 1.010 1.400 1.740 ;
        RECT  0.120 1.500 1.400 1.740 ;
        RECT  1.890 1.010 2.130 1.990 ;
        RECT  1.890 1.750 2.960 1.990 ;
        RECT  0.120 1.500 0.830 2.100 ;
        RECT  2.720 1.750 2.960 2.490 ;
        RECT  0.120 1.500 0.360 3.540 ;
        RECT  0.230 3.300 0.510 3.850 ;
        RECT  3.050 0.980 3.630 1.460 ;
        RECT  3.190 0.980 3.630 3.230 ;
        RECT  3.190 1.850 4.650 2.250 ;
        RECT  3.190 1.850 3.640 3.230 ;
        RECT  2.890 2.730 3.270 4.610 ;
        RECT  2.840 3.920 3.270 4.610 ;
    END
END nr03da

MACRO nr03d7
    CLASS CORE ;
    FOREIGN nr03d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.610 2.350 1.060 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.467  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.690 1.620 4.140 ;
        RECT  1.350 1.980 1.620 4.140 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.467  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.040 3.080 2.740 3.600 ;
        RECT  2.040 2.260 2.280 3.600 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.451  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.480 1.340 7.530 1.580 ;
        RECT  6.470 1.340 6.870 2.940 ;
        RECT  5.430 2.640 6.870 2.880 ;
        RECT  6.220 1.340 6.870 2.880 ;
        RECT  5.430 2.640 5.670 4.310 ;
        RECT  4.110 3.420 5.670 3.660 ;
        RECT  4.110 3.420 4.350 4.590 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  7.250 4.620 7.650 5.600 ;
        RECT  5.910 3.230 6.310 5.600 ;
        RECT  4.790 4.620 5.190 5.600 ;
        RECT  3.460 3.470 3.870 5.600 ;
        RECT  2.020 4.620 2.420 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.340 0.000 6.740 0.980 ;
        RECT  5.040 0.000 5.440 0.980 ;
        RECT  3.740 0.000 4.140 0.980 ;
        RECT  2.390 0.000 2.630 1.330 ;
        RECT  0.270 1.010 0.830 1.260 ;
        RECT  0.270 0.000 0.510 1.260 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.160 1.010 2.130 1.250 ;
        RECT  1.160 1.010 1.400 1.740 ;
        RECT  0.120 1.500 1.400 1.740 ;
        RECT  1.890 1.010 2.130 1.990 ;
        RECT  1.890 1.750 2.960 1.990 ;
        RECT  0.120 1.500 0.830 2.100 ;
        RECT  2.720 1.750 2.960 2.490 ;
        RECT  0.120 1.500 0.360 3.540 ;
        RECT  0.230 3.300 0.510 3.850 ;
        RECT  3.050 0.980 3.440 1.380 ;
        RECT  3.200 1.990 5.980 2.390 ;
        RECT  3.200 0.980 3.440 2.970 ;
        RECT  2.980 2.730 3.220 4.160 ;
        RECT  2.840 3.920 3.080 4.610 ;
    END
END nr03d7

MACRO nr03d4
    CLASS CORE ;
    FOREIGN nr03d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.700 1.060 4.140 ;
        RECT  0.710 2.520 0.950 4.140 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.190 2.520 1.720 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.527  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.000 2.520 2.740 3.020 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.857  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.250 3.130 6.010 3.370 ;
        RECT  4.230 1.600 6.010 1.840 ;
        RECT  5.100 1.600 5.540 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.930 4.570 5.330 5.600 ;
        RECT  3.510 4.570 3.910 5.600 ;
        RECT  2.110 4.230 2.350 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.000 0.000 5.400 1.010 ;
        RECT  3.550 0.000 3.950 1.060 ;
        RECT  2.270 0.000 2.510 1.510 ;
        RECT  0.880 0.000 1.120 1.510 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.770 0.550 2.090 ;
        RECT  0.150 1.850 3.410 2.090 ;
        RECT  0.150 1.770 0.470 2.170 ;
        RECT  0.230 1.770 0.470 3.450 ;
        RECT  2.890 1.320 3.890 1.560 ;
        RECT  3.650 2.320 4.380 2.560 ;
        RECT  3.650 1.320 3.890 3.500 ;
        RECT  2.870 3.260 3.890 3.500 ;
    END
END nr03d4

MACRO nr03d2
    CLASS CORE ;
    FOREIGN nr03d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.700 1.060 4.140 ;
        RECT  0.710 2.520 0.950 4.140 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.190 2.520 1.720 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.527  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.080 3.140 2.740 3.580 ;
        RECT  2.080 2.520 2.320 3.580 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.248  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.310 3.140 4.980 3.580 ;
        RECT  4.740 1.850 4.980 3.580 ;
        RECT  4.370 1.850 4.980 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  5.100 4.070 5.340 5.600 ;
        RECT  3.770 4.070 4.010 5.600 ;
        RECT  2.110 4.230 2.350 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  5.050 0.000 5.450 0.890 ;
        RECT  3.590 0.000 4.030 0.890 ;
        RECT  2.270 0.000 2.510 1.510 ;
        RECT  0.880 0.000 1.120 1.510 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.770 0.550 2.090 ;
        RECT  0.150 1.850 2.770 2.090 ;
        RECT  2.530 1.850 2.770 2.400 ;
        RECT  0.150 1.770 0.470 2.170 ;
        RECT  2.530 2.160 3.450 2.400 ;
        RECT  0.230 1.770 0.470 3.450 ;
        RECT  2.970 1.470 3.930 1.710 ;
        RECT  3.690 2.380 4.460 2.620 ;
        RECT  3.690 1.470 3.930 3.370 ;
        RECT  3.090 3.130 3.930 3.370 ;
        RECT  3.090 3.130 3.330 3.690 ;
    END
END nr03d2

MACRO nr03d1
    CLASS CORE ;
    FOREIGN nr03d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.300 2.180 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.700 1.600 4.150 ;
        RECT  1.230 2.520 1.470 4.150 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.500 3.020 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.733  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.200 1.820 2.680 2.060 ;
        RECT  2.300 1.460 2.680 2.060 ;
        RECT  0.200 3.260 0.980 3.500 ;
        RECT  0.740 1.820 0.980 3.500 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  1.890 4.710 2.320 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  2.250 0.000 2.650 0.890 ;
        RECT  0.800 0.000 1.040 1.420 ;
        END
    END VSS
END nr03d1

MACRO nr03d0
    CLASS CORE ;
    FOREIGN nr03d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.238  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.180 3.580 ;
        RECT  1.840 2.580 2.080 3.580 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.238  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 2.020 1.620 2.460 ;
        RECT  1.160 2.020 1.400 2.980 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.238  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.180 0.800 2.500 ;
        RECT  0.120 2.180 0.500 3.020 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.942  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.230 3.820 2.680 4.060 ;
        RECT  2.420 1.540 2.680 4.060 ;
        RECT  2.300 1.540 2.680 2.460 ;
        RECT  0.150 1.540 2.680 1.780 ;
        RECT  0.230 3.500 0.470 4.060 ;
        RECT  0.150 1.540 0.470 1.940 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  2.060 4.710 2.490 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  2.200 0.000 2.600 0.890 ;
        RECT  0.570 0.000 0.970 0.890 ;
        END
    END VSS
END nr03d0

MACRO nr02da
    CLASS CORE ;
    FOREIGN nr02da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.700 2.660 2.460 ;
        RECT  1.290 1.700 2.660 2.100 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.471  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.890 0.550 2.530 ;
        RECT  0.120 1.890 0.500 3.020 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.659  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.510 1.390 8.840 2.940 ;
        RECT  8.230 1.390 8.730 3.450 ;
        RECT  7.500 1.310 7.900 2.940 ;
        RECT  7.010 1.390 7.580 4.620 ;
        RECT  6.020 1.310 6.420 2.940 ;
        RECT  5.700 1.390 6.200 4.340 ;
        RECT  3.540 2.740 6.200 3.190 ;
        RECT  4.580 1.390 5.090 4.550 ;
        RECT  4.510 1.150 4.940 3.240 ;
        RECT  3.540 2.740 5.090 3.240 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.920 3.720 8.160 5.600 ;
        RECT  6.520 3.260 6.760 5.600 ;
        RECT  5.320 4.620 5.720 5.600 ;
        RECT  4.100 3.470 4.340 5.600 ;
        RECT  2.800 4.450 3.040 5.600 ;
        RECT  1.560 2.630 1.800 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  8.240 0.000 8.640 0.980 ;
        RECT  6.760 0.000 7.160 1.010 ;
        RECT  5.280 0.000 5.680 1.090 ;
        RECT  3.800 0.000 4.200 0.980 ;
        RECT  1.730 0.000 2.130 0.890 ;
        RECT  0.300 0.000 0.540 1.430 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.800 1.140 2.660 1.380 ;
        RECT  0.800 1.110 1.510 1.430 ;
        RECT  0.800 1.110 1.040 4.540 ;
        RECT  0.150 4.300 1.040 4.540 ;
        RECT  2.890 0.980 3.300 3.500 ;
        RECT  2.890 2.060 4.280 2.510 ;
        RECT  2.890 2.060 3.310 3.500 ;
        RECT  2.190 3.000 3.310 3.500 ;
    END
END nr02da

MACRO nr02d7
    CLASS CORE ;
    FOREIGN nr02d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.700 2.740 2.460 ;
        RECT  1.290 1.700 2.740 2.100 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.471  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.890 0.550 2.530 ;
        RECT  0.120 1.890 0.500 3.020 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.669  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.540 2.680 7.160 3.080 ;
        RECT  6.780 1.370 7.160 3.080 ;
        RECT  4.480 1.370 7.160 1.770 ;
        RECT  5.950 4.220 6.520 4.620 ;
        RECT  5.950 2.680 6.190 4.620 ;
        RECT  4.870 2.680 5.110 4.450 ;
        RECT  3.540 2.680 3.780 4.420 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.810 3.550 7.050 5.600 ;
        RECT  5.460 3.380 5.700 5.600 ;
        RECT  4.130 3.330 4.370 5.600 ;
        RECT  2.800 3.930 3.040 5.600 ;
        RECT  1.560 2.630 1.800 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.570 0.000 6.970 1.010 ;
        RECT  5.220 0.000 5.620 1.090 ;
        RECT  3.790 0.000 4.190 1.070 ;
        RECT  1.730 0.000 2.130 0.890 ;
        RECT  0.300 0.000 0.540 1.430 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.800 1.140 2.660 1.380 ;
        RECT  0.800 1.030 1.510 1.430 ;
        RECT  0.800 1.030 1.040 4.540 ;
        RECT  0.150 4.300 1.040 4.540 ;
        RECT  2.900 0.980 3.300 1.390 ;
        RECT  2.980 2.010 6.340 2.410 ;
        RECT  2.980 0.980 3.220 3.500 ;
        RECT  2.190 3.260 3.220 3.500 ;
    END
END nr02d7

MACRO nr02d4
    CLASS CORE ;
    FOREIGN nr02d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.450 3.020 ;
        RECT  1.210 2.180 1.450 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.100 0.830 2.340 ;
        RECT  0.120 1.460 0.500 2.340 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.143  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.740 3.130 5.440 3.370 ;
        RECT  3.740 1.710 5.440 1.950 ;
        RECT  4.540 1.710 4.980 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.270 4.620 4.670 5.600 ;
        RECT  2.970 4.620 3.370 5.600 ;
        RECT  1.410 4.710 1.810 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.480 0.000 4.880 0.980 ;
        RECT  3.150 0.000 3.550 0.910 ;
        RECT  1.710 0.000 2.110 0.890 ;
        RECT  0.150 0.000 0.550 0.900 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.920 1.570 2.010 1.810 ;
        RECT  1.770 2.260 2.780 2.500 ;
        RECT  1.770 1.570 2.010 3.500 ;
        RECT  0.180 3.260 2.010 3.500 ;
        RECT  2.350 1.730 3.260 1.970 ;
        RECT  3.020 2.260 3.860 2.500 ;
        RECT  3.020 1.730 3.260 3.370 ;
        RECT  2.350 3.130 3.260 3.370 ;
    END
END nr02d4

MACRO nr02d2
    CLASS CORE ;
    FOREIGN nr02d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.002  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.580 2.050 2.840 ;
        RECT  1.180 2.580 1.620 3.040 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.723  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.380 0.870 2.620 ;
        RECT  0.120 2.380 0.500 3.020 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.775  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.550 3.280 2.740 3.520 ;
        RECT  2.300 1.660 2.740 3.520 ;
        RECT  0.720 1.770 2.740 2.010 ;
        RECT  2.070 1.660 2.740 2.010 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.870 4.160 3.110 5.600 ;
        RECT  0.610 4.160 0.850 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.890 0.000 3.130 1.420 ;
        RECT  1.540 0.000 1.780 1.420 ;
        RECT  0.230 0.000 0.470 1.420 ;
        END
    END VSS
END nr02d2

MACRO nr02d1
    CLASS CORE ;
    FOREIGN nr02d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.580 1.620 3.020 ;
        RECT  1.180 2.020 1.440 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.100 0.820 2.340 ;
        RECT  0.120 2.100 0.500 3.020 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.390  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.170 3.260 2.120 3.500 ;
        RECT  1.860 1.220 2.120 3.500 ;
        RECT  1.740 1.220 2.120 1.900 ;
        RECT  0.990 1.220 2.120 1.460 ;
        RECT  0.990 1.220 1.230 1.780 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.240 5.600 ;
        RECT  1.670 4.710 2.090 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.240 0.740 ;
        RECT  1.680 0.000 2.090 0.890 ;
        RECT  0.230 0.000 0.470 1.420 ;
        END
    END VSS
END nr02d1

MACRO nr02d0
    CLASS CORE ;
    FOREIGN nr02d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.100 0.820 2.340 ;
        RECT  0.120 2.100 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.580 1.620 3.020 ;
        RECT  1.180 2.020 1.440 3.020 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.705  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.170 3.260 2.120 3.500 ;
        RECT  1.860 1.230 2.120 3.500 ;
        RECT  1.740 1.230 2.120 1.900 ;
        RECT  0.990 1.230 2.120 1.470 ;
        RECT  0.990 1.230 1.230 1.780 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.240 5.600 ;
        RECT  1.400 4.710 1.800 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.240 0.740 ;
        RECT  1.680 0.000 2.080 0.990 ;
        RECT  0.230 0.000 0.470 1.720 ;
        END
    END VSS
END nr02d0

MACRO nd23d4
    CLASS CORE ;
    FOREIGN nd23d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.301  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.020 3.210 2.620 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.301  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.470 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.290 0.710 2.610 ;
        RECT  0.120 2.290 0.500 3.020 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.837  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.150 3.190 5.910 3.430 ;
        RECT  4.150 1.600 5.910 1.840 ;
        RECT  5.100 1.600 5.540 3.430 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.830 4.570 5.230 5.600 ;
        RECT  3.380 4.570 3.780 5.600 ;
        RECT  0.300 3.270 0.540 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.920 0.000 5.320 0.890 ;
        RECT  3.500 0.000 3.930 0.890 ;
        RECT  1.790 0.000 2.190 0.890 ;
        RECT  0.300 0.000 0.550 2.050 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.070 2.490 1.660 2.730 ;
        RECT  1.070 1.740 1.310 3.470 ;
        RECT  1.020 0.980 1.340 1.370 ;
        RECT  2.560 0.980 2.960 1.370 ;
        RECT  1.020 1.130 3.690 1.370 ;
        RECT  3.450 2.320 4.300 2.560 ;
        RECT  3.450 1.130 3.690 4.170 ;
        RECT  1.110 3.930 3.690 4.170 ;
    END
END nd23d4

MACRO nd23d2
    CLASS CORE ;
    FOREIGN nd23d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.301  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.020 3.210 2.620 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.301  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.470 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.290 0.710 2.610 ;
        RECT  0.120 2.290 0.500 3.020 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 3.140 4.560 3.940 ;
        RECT  4.320 1.450 4.560 3.940 ;
        RECT  4.100 1.450 4.560 1.780 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.840 4.530 5.240 5.600 ;
        RECT  3.360 4.530 3.760 5.600 ;
        RECT  0.300 3.270 0.540 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.920 0.000 5.160 1.280 ;
        RECT  3.330 0.000 3.730 0.890 ;
        RECT  1.790 0.000 2.190 0.890 ;
        RECT  0.300 0.000 0.540 2.050 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.070 2.490 1.660 2.730 ;
        RECT  1.070 1.740 1.310 3.470 ;
        RECT  1.020 0.980 1.340 1.370 ;
        RECT  2.560 0.980 2.960 1.370 ;
        RECT  1.020 1.130 3.690 1.370 ;
        RECT  3.450 2.380 4.080 2.620 ;
        RECT  3.450 1.130 3.690 4.170 ;
        RECT  1.110 3.930 3.690 4.170 ;
    END
END nd23d2

MACRO nd23d1
    CLASS CORE ;
    FOREIGN nd23d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.106  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.700 1.670 4.150 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.500 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.910 2.020 4.420 2.790 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.783  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.210 3.130 3.990 3.370 ;
        RECT  2.860 3.130 3.300 3.580 ;
        RECT  2.740 1.850 2.980 3.370 ;
        RECT  2.210 1.850 2.980 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.270 4.130 4.510 5.600 ;
        RECT  2.900 4.130 3.140 5.600 ;
        RECT  0.640 4.510 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.200 0.000 4.440 1.480 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 2.470 2.500 2.710 ;
        RECT  1.590 1.770 1.830 3.460 ;
        RECT  0.740 1.290 3.460 1.530 ;
        RECT  0.150 1.730 0.980 1.970 ;
        RECT  3.220 1.290 3.460 2.800 ;
        RECT  0.740 1.290 0.980 3.500 ;
        RECT  0.150 3.260 0.980 3.500 ;
    END
END nd23d1

MACRO nd13d4
    CLASS CORE ;
    FOREIGN nd13d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.340 0.800 2.580 ;
        RECT  0.120 2.340 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.500 2.250 2.940 2.650 ;
        RECT  2.500 1.460 2.740 2.650 ;
        RECT  2.300 1.460 2.740 1.900 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.150 2.180 3.020 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.020 3.130 6.720 3.370 ;
        RECT  4.950 1.850 6.720 2.090 ;
        RECT  5.660 1.850 6.100 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  5.630 4.570 6.040 5.600 ;
        RECT  4.280 4.570 4.680 5.600 ;
        RECT  2.190 4.570 2.590 5.600 ;
        RECT  0.870 4.360 1.110 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  5.640 0.000 6.040 0.890 ;
        RECT  4.220 0.000 4.620 0.890 ;
        RECT  0.750 0.000 1.150 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.690 1.280 1.930 ;
        RECT  1.040 2.160 1.480 2.550 ;
        RECT  1.040 1.690 1.280 3.500 ;
        RECT  0.150 3.260 1.280 3.500 ;
        RECT  2.980 1.460 3.220 2.010 ;
        RECT  3.180 2.450 4.210 2.690 ;
        RECT  3.180 1.770 3.420 3.500 ;
        RECT  1.570 3.260 3.420 3.500 ;
        RECT  3.680 1.600 4.690 1.840 ;
        RECT  3.680 1.600 3.920 2.160 ;
        RECT  4.450 2.380 5.050 2.620 ;
        RECT  3.680 3.050 3.920 3.640 ;
        RECT  4.450 1.600 4.690 3.640 ;
        RECT  3.680 3.400 4.690 3.640 ;
    END
END nd13d4

MACRO nd13d2
    CLASS CORE ;
    FOREIGN nd13d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.770 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.767  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.680 2.580 2.180 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.994  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.600 2.580 3.300 3.020 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.670  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.640 3.270 4.980 3.510 ;
        RECT  4.740 1.440 4.980 3.510 ;
        RECT  4.540 1.440 4.980 2.460 ;
        RECT  2.950 1.440 4.980 1.680 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  5.110 4.300 5.350 5.600 ;
        RECT  3.780 4.300 4.020 5.600 ;
        RECT  2.480 4.300 2.720 5.600 ;
        RECT  1.130 4.270 1.370 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.660 0.000 5.060 0.890 ;
        RECT  1.150 0.000 1.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.280 1.500 1.020 1.740 ;
        RECT  0.780 2.030 4.300 2.270 ;
        RECT  4.060 2.030 4.300 3.030 ;
        RECT  0.780 1.500 1.020 3.480 ;
        RECT  0.280 3.240 1.020 3.480 ;
    END
END nd13d2

MACRO nd13d1
    CLASS CORE ;
    FOREIGN nd13d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.340 0.800 2.580 ;
        RECT  0.120 2.340 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.500 2.250 2.940 2.650 ;
        RECT  2.500 1.460 2.740 2.650 ;
        RECT  2.300 1.460 2.740 1.900 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.150 2.180 3.020 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.769  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 3.140 3.420 3.580 ;
        RECT  3.180 1.770 3.420 3.580 ;
        RECT  2.980 1.460 3.220 2.010 ;
        RECT  1.570 3.260 3.420 3.500 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  2.270 4.370 2.510 5.600 ;
        RECT  0.870 4.360 1.110 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  0.750 0.000 1.150 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.690 1.280 1.930 ;
        RECT  1.040 2.160 1.480 2.550 ;
        RECT  1.040 1.690 1.280 3.500 ;
        RECT  0.150 3.260 1.280 3.500 ;
    END
END nd13d1

MACRO nd12d4
    CLASS CORE ;
    FOREIGN nd12d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.160 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.160 2.180 3.020 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.310 3.130 6.010 3.370 ;
        RECT  4.240 1.850 6.010 2.090 ;
        RECT  5.100 1.850 5.540 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.920 4.570 5.330 5.600 ;
        RECT  3.570 4.570 3.970 5.600 ;
        RECT  2.270 4.060 2.510 5.600 ;
        RECT  0.860 4.710 1.260 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.930 0.000 5.330 0.890 ;
        RECT  3.510 0.000 3.910 0.890 ;
        RECT  0.960 0.000 1.360 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.680 1.430 1.920 ;
        RECT  1.190 1.680 1.430 3.020 ;
        RECT  0.740 2.780 1.430 3.020 ;
        RECT  0.740 2.780 0.980 3.500 ;
        RECT  0.150 3.260 0.980 3.500 ;
        RECT  2.190 1.600 2.660 1.920 ;
        RECT  2.420 2.450 3.500 2.690 ;
        RECT  2.420 1.600 2.660 3.500 ;
        RECT  1.600 3.260 2.660 3.500 ;
        RECT  2.970 1.600 3.980 1.840 ;
        RECT  2.970 1.600 3.210 2.170 ;
        RECT  3.740 2.380 4.340 2.620 ;
        RECT  2.970 3.050 3.210 3.600 ;
        RECT  3.740 1.600 3.980 3.600 ;
        RECT  2.970 3.360 3.980 3.600 ;
    END
END nd12d4

MACRO nd12d2
    CLASS CORE ;
    FOREIGN nd12d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.925  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.120 2.020 2.740 2.700 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.128  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 3.140 3.520 3.580 ;
        RECT  2.980 3.050 3.520 3.580 ;
        RECT  2.980 1.490 3.220 3.580 ;
        RECT  2.380 1.490 3.220 1.740 ;
        RECT  1.640 3.140 3.520 3.380 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.760 4.160 4.000 5.600 ;
        RECT  2.460 4.160 2.700 5.600 ;
        RECT  0.870 4.160 1.110 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.660 0.000 3.900 1.560 ;
        RECT  1.130 0.000 1.370 1.540 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.210 1.780 0.980 2.020 ;
        RECT  0.740 2.380 1.540 2.620 ;
        RECT  0.740 1.780 0.980 3.500 ;
        RECT  0.210 3.260 0.980 3.500 ;
    END
END nd12d2

MACRO nd12d1
    CLASS CORE ;
    FOREIGN nd12d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.309  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.140 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.200 3.020 ;
        RECT  1.960 2.140 2.200 3.020 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.660 3.260 2.680 3.500 ;
        RECT  2.440 1.460 2.680 3.500 ;
        RECT  2.250 1.460 2.680 1.900 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  2.330 4.080 2.570 5.600 ;
        RECT  1.030 4.080 1.270 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  0.920 0.000 1.320 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.660 1.490 1.900 ;
        RECT  1.250 1.660 1.490 3.020 ;
        RECT  0.740 2.780 1.490 3.020 ;
        RECT  0.740 2.780 0.980 3.500 ;
        RECT  0.160 3.260 0.980 3.500 ;
    END
END nd12d1

MACRO nd12d0
    CLASS CORE ;
    FOREIGN nd12d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.340 0.810 2.580 ;
        RECT  0.120 2.340 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.200 3.020 ;
        RECT  1.960 2.130 2.200 3.020 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.582  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.530 3.260 2.680 3.500 ;
        RECT  2.440 1.140 2.680 3.500 ;
        RECT  2.300 1.140 2.680 1.900 ;
        RECT  2.130 1.140 2.680 1.460 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  2.130 4.710 2.530 5.600 ;
        RECT  0.570 4.710 0.970 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  0.990 0.000 1.230 1.540 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.200 0.470 2.100 ;
        RECT  0.230 1.860 1.290 2.100 ;
        RECT  1.050 2.000 1.580 2.400 ;
        RECT  1.050 1.860 1.290 3.500 ;
        RECT  0.170 3.260 1.290 3.500 ;
    END
END nd12d0

MACRO nd04da
    CLASS CORE ;
    FOREIGN nd04da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.353  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.250 3.580 ;
        RECT  1.010 2.620 1.250 3.580 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.440 2.520 3.380 3.040 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.660 1.990 2.180 3.110 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.353  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.970 0.640 2.800 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.045  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.800 3.930 9.470 4.330 ;
        RECT  9.070 1.170 9.470 4.330 ;
        RECT  5.030 2.590 9.470 4.330 ;
        RECT  5.970 1.250 9.470 4.330 ;
        RECT  7.560 1.170 7.960 4.330 ;
        RECT  4.590 1.210 6.470 1.710 ;
        RECT  6.070 1.170 6.470 4.330 ;
        RECT  4.590 1.000 5.040 1.710 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  9.460 4.600 9.900 5.600 ;
        RECT  8.130 4.610 8.540 5.600 ;
        RECT  6.840 4.620 7.240 5.600 ;
        RECT  5.540 4.620 5.940 5.600 ;
        RECT  4.170 4.700 4.570 5.600 ;
        RECT  2.870 4.650 3.270 5.600 ;
        RECT  1.290 4.710 1.690 5.600 ;
        RECT  0.150 4.710 0.590 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  8.300 0.000 8.700 0.980 ;
        RECT  6.810 0.000 7.210 0.980 ;
        RECT  5.330 0.000 5.730 0.980 ;
        RECT  3.850 0.000 4.250 0.980 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.250 1.490 2.850 1.730 ;
        RECT  2.610 1.490 2.850 2.240 ;
        RECT  2.610 2.000 3.860 2.240 ;
        RECT  3.620 2.000 3.860 3.590 ;
        RECT  1.660 3.350 3.860 3.590 ;
        RECT  1.660 3.350 1.900 4.080 ;
        RECT  0.710 3.840 1.900 4.080 ;
        RECT  3.120 1.130 3.520 1.750 ;
        RECT  3.120 1.350 4.350 1.750 ;
        RECT  4.100 1.350 4.350 4.230 ;
        RECT  4.100 1.940 5.740 2.340 ;
        RECT  4.100 1.940 4.500 4.230 ;
        RECT  3.460 3.830 4.500 4.230 ;
    END
END nd04da

MACRO nd04d7
    CLASS CORE ;
    FOREIGN nd04d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.990 2.180 3.110 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.970 0.640 2.800 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.400 3.580 ;
        RECT  1.050 2.620 1.400 3.580 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.440 2.480 3.380 3.040 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.982  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.920 1.150 8.650 1.550 ;
        RECT  4.790 3.920 8.340 4.320 ;
        RECT  7.900 1.150 8.340 4.320 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  8.230 4.620 8.630 5.600 ;
        RECT  6.840 4.620 7.240 5.600 ;
        RECT  5.540 4.620 5.940 5.600 ;
        RECT  4.170 4.700 4.570 5.600 ;
        RECT  2.870 4.650 3.270 5.600 ;
        RECT  1.010 4.600 1.410 5.600 ;
        RECT  0.150 4.710 0.590 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.330 0.000 7.730 0.890 ;
        RECT  5.690 0.000 6.090 0.890 ;
        RECT  4.180 0.000 4.580 0.980 ;
        RECT  2.450 0.000 2.850 0.950 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.490 2.760 1.730 ;
        RECT  2.520 1.490 2.760 2.230 ;
        RECT  2.520 1.990 3.980 2.230 ;
        RECT  3.740 1.990 3.980 3.590 ;
        RECT  1.660 3.350 3.980 3.590 ;
        RECT  1.660 3.350 1.900 4.080 ;
        RECT  0.710 3.840 1.900 4.080 ;
        RECT  3.300 1.010 3.540 1.730 ;
        RECT  3.300 1.490 4.460 1.730 ;
        RECT  4.220 1.810 7.150 2.210 ;
        RECT  4.220 1.490 4.460 4.230 ;
        RECT  3.460 3.990 4.460 4.230 ;
    END
END nd04d7

MACRO nd04d4
    CLASS CORE ;
    FOREIGN nd04d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.460 1.620 1.900 ;
        RECT  1.160 1.460 1.400 2.640 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.460 2.760 2.920 ;
        RECT  2.300 1.460 2.760 1.900 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.240 2.180 3.020 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.230 0.500 3.020 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.870 3.130 6.570 3.370 ;
        RECT  4.800 1.850 6.570 2.090 ;
        RECT  5.660 1.850 6.100 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.490 4.570 5.890 5.600 ;
        RECT  4.130 4.570 4.530 5.600 ;
        RECT  2.680 4.710 3.080 5.600 ;
        RECT  1.590 4.390 1.830 5.600 ;
        RECT  0.240 4.710 0.640 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.570 0.000 5.810 1.330 ;
        RECT  4.150 0.000 4.390 1.330 ;
        RECT  0.230 0.000 0.470 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.720 0.980 3.280 1.220 ;
        RECT  3.030 0.980 3.280 2.690 ;
        RECT  3.030 2.450 4.060 2.690 ;
        RECT  3.030 0.980 3.270 3.500 ;
        RECT  0.740 3.260 3.270 3.500 ;
        RECT  3.530 1.610 4.540 1.850 ;
        RECT  3.530 1.610 3.770 2.170 ;
        RECT  4.300 2.380 4.900 2.620 ;
        RECT  3.530 3.050 3.770 3.600 ;
        RECT  4.300 1.610 4.540 3.600 ;
        RECT  3.530 3.360 4.540 3.600 ;
    END
END nd04d4

MACRO nd04d2
    CLASS CORE ;
    FOREIGN nd04d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.460 1.620 1.900 ;
        RECT  1.150 1.460 1.400 2.640 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.500 1.460 2.790 2.920 ;
        RECT  2.300 1.460 2.790 1.900 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.240 2.180 3.020 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.230 0.500 3.020 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.251  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.790 3.130 5.540 3.370 ;
        RECT  5.100 1.850 5.540 3.370 ;
        RECT  4.790 1.850 5.540 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.490 4.710 5.890 5.600 ;
        RECT  4.130 4.710 4.530 5.600 ;
        RECT  2.680 4.710 3.080 5.600 ;
        RECT  1.590 4.390 1.830 5.600 ;
        RECT  0.240 4.710 0.640 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.570 0.000 5.810 1.600 ;
        RECT  4.150 0.000 4.390 1.370 ;
        RECT  0.230 0.000 0.470 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.720 0.980 3.270 1.220 ;
        RECT  3.030 2.450 4.060 2.690 ;
        RECT  3.030 0.980 3.270 3.500 ;
        RECT  0.740 3.260 3.270 3.500 ;
        RECT  3.520 1.610 4.540 1.850 ;
        RECT  3.520 1.610 3.760 2.170 ;
        RECT  4.300 2.380 4.860 2.620 ;
        RECT  3.530 3.050 3.770 3.600 ;
        RECT  4.300 1.610 4.540 3.600 ;
        RECT  3.530 3.360 4.540 3.600 ;
    END
END nd04d2

MACRO nd04d1
    CLASS CORE ;
    FOREIGN nd04d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.460 1.460 2.640 ;
        RECT  0.620 1.460 1.460 1.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.240 2.690 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.820 2.140 2.640 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.320 0.500 3.020 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.853  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.540 3.160 1.780 ;
        RECT  2.220 3.140 2.740 3.580 ;
        RECT  0.740 3.130 2.620 3.370 ;
        RECT  2.380 1.540 2.620 3.580 ;
        RECT  2.220 3.050 2.620 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.740 4.710 3.140 5.600 ;
        RECT  1.610 4.300 1.850 5.600 ;
        RECT  0.240 4.710 0.640 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  0.180 0.000 0.580 0.890 ;
        END
    END VSS
END nd04d1

MACRO nd04d0
    CLASS CORE ;
    FOREIGN nd04d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.580 1.620 3.020 ;
        RECT  1.180 2.090 1.540 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.240 2.730 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.460 2.140 2.490 ;
        RECT  1.740 1.460 2.140 1.900 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.390 0.500 3.580 ;
        END
    END A4
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.000  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.540 3.120 1.780 ;
        RECT  2.220 3.140 2.740 3.580 ;
        RECT  2.380 1.540 2.620 3.580 ;
        RECT  0.740 3.260 2.740 3.500 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.890 4.300 3.130 5.600 ;
        RECT  1.590 4.300 1.830 5.600 ;
        RECT  0.230 4.300 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
END nd04d0

MACRO nd03da
    CLASS CORE ;
    FOREIGN nd03da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.340 0.800 2.740 ;
        RECT  0.120 2.020 0.500 2.740 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.040 2.020 1.540 2.630 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 2.020 2.240 2.630 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.546  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.780 1.220 9.180 1.620 ;
        RECT  5.180 1.270 9.100 2.460 ;
        RECT  8.560 1.240 9.180 1.620 ;
        RECT  4.240 2.870 8.540 4.020 ;
        RECT  5.180 1.270 8.540 4.020 ;
        RECT  4.240 1.240 7.800 1.740 ;
        RECT  7.300 1.210 7.700 4.020 ;
        RECT  5.820 1.210 6.220 4.020 ;
        RECT  4.340 1.220 4.740 1.740 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  8.860 3.050 9.260 5.600 ;
        RECT  7.580 4.620 7.980 5.600 ;
        RECT  6.280 4.620 6.680 5.600 ;
        RECT  4.980 4.620 5.380 5.600 ;
        RECT  3.670 4.620 4.070 5.600 ;
        RECT  2.150 3.350 2.550 5.600 ;
        RECT  0.570 4.710 0.970 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.040 0.000 8.440 1.040 ;
        RECT  6.560 0.000 6.960 1.010 ;
        RECT  5.080 0.000 5.480 1.010 ;
        RECT  3.590 0.000 4.000 0.990 ;
        RECT  2.140 0.000 2.540 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.170 1.290 1.510 1.530 ;
        RECT  1.270 1.290 1.510 1.780 ;
        RECT  1.270 1.540 2.670 1.780 ;
        RECT  2.480 1.590 2.720 2.030 ;
        RECT  2.600 1.790 2.840 3.110 ;
        RECT  1.490 2.870 2.840 3.110 ;
        RECT  0.150 3.210 1.730 3.460 ;
        RECT  1.490 2.870 1.730 4.350 ;
        RECT  2.890 0.980 3.360 1.380 ;
        RECT  3.080 0.980 3.360 3.900 ;
        RECT  3.080 1.970 4.950 2.380 ;
        RECT  3.080 1.970 3.480 3.900 ;
        RECT  2.900 3.500 3.480 3.900 ;
    END
END nd03da

MACRO nd03d7
    CLASS CORE ;
    FOREIGN nd03d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.340 0.720 2.740 ;
        RECT  0.120 2.010 0.500 2.740 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.100 1.950 1.540 2.610 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 2.020 2.200 2.630 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.738  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.650 2.500 7.690 2.810 ;
        RECT  7.290 1.220 7.690 2.810 ;
        RECT  4.330 1.300 7.690 1.540 ;
        RECT  6.650 2.500 7.050 4.150 ;
        RECT  4.040 3.360 7.050 3.760 ;
        RECT  6.210 3.140 7.050 3.760 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  7.290 3.050 7.690 5.600 ;
        RECT  6.080 4.620 6.480 5.600 ;
        RECT  4.780 4.620 5.180 5.600 ;
        RECT  3.550 4.280 3.790 5.600 ;
        RECT  2.230 3.350 2.470 5.600 ;
        RECT  2.070 3.350 2.470 3.750 ;
        RECT  0.590 4.710 0.990 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.550 0.000 6.950 1.050 ;
        RECT  5.070 0.000 5.470 1.050 ;
        RECT  3.670 0.000 3.910 1.060 ;
        RECT  2.110 0.000 2.540 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.170 1.210 0.570 1.700 ;
        RECT  0.170 1.460 1.900 1.700 ;
        RECT  1.720 1.540 2.840 1.780 ;
        RECT  2.600 1.540 2.840 3.110 ;
        RECT  1.420 2.870 2.840 3.110 ;
        RECT  1.420 2.870 1.660 3.460 ;
        RECT  0.150 3.210 1.660 3.460 ;
        RECT  1.190 3.210 1.430 4.350 ;
        RECT  1.190 4.110 1.880 4.350 ;
        RECT  2.880 1.060 3.430 1.300 ;
        RECT  3.190 1.860 7.000 2.260 ;
        RECT  3.190 1.060 3.430 4.010 ;
        RECT  3.070 3.770 3.310 4.590 ;
        RECT  2.750 4.350 3.310 4.590 ;
    END
END nd03d7

MACRO nd03d4
    CLASS CORE ;
    FOREIGN nd03d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.100 0.810 2.340 ;
        RECT  0.120 2.100 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 1.900 ;
        RECT  1.180 1.460 1.420 2.380 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.180 3.020 ;
        RECT  1.900 1.980 2.180 3.020 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.230 3.130 5.940 3.370 ;
        RECT  4.170 1.850 5.940 2.090 ;
        RECT  4.540 1.850 4.980 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.860 4.570 5.260 5.600 ;
        RECT  3.500 4.570 3.900 5.600 ;
        RECT  2.080 4.430 2.480 5.600 ;
        RECT  1.360 4.400 1.600 5.600 ;
        RECT  0.590 3.250 0.830 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.860 0.000 5.260 0.890 ;
        RECT  3.440 0.000 3.840 0.890 ;
        RECT  0.160 0.000 0.570 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.080 1.500 2.660 1.740 ;
        RECT  2.420 2.450 3.430 2.690 ;
        RECT  2.420 1.500 2.660 3.550 ;
        RECT  1.350 3.310 2.660 3.550 ;
        RECT  2.900 1.610 3.910 1.850 ;
        RECT  2.900 1.610 3.140 2.170 ;
        RECT  3.670 2.380 4.270 2.620 ;
        RECT  2.900 3.050 3.140 3.600 ;
        RECT  3.670 1.610 3.910 3.600 ;
        RECT  2.900 3.360 3.910 3.600 ;
    END
END nd03d4

MACRO nd03d2
    CLASS CORE ;
    FOREIGN nd03d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.806  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.410 3.860 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.982  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.540 3.080 2.460 ;
        RECT  0.120 1.540 3.080 1.780 ;
        RECT  0.120 1.540 0.500 2.910 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.983  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.220 2.080 2.460 ;
        RECT  1.180 2.020 1.620 2.460 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.995  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.720 3.260 4.920 3.500 ;
        RECT  4.540 1.830 4.920 3.500 ;
        RECT  3.320 1.830 4.920 2.070 ;
        RECT  3.320 1.060 3.560 2.070 ;
        RECT  1.810 1.060 3.560 1.300 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.180 4.030 4.420 5.600 ;
        RECT  2.840 4.210 3.080 5.600 ;
        RECT  1.540 4.210 1.780 5.600 ;
        RECT  0.230 4.210 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.820 0.000 4.060 1.470 ;
        RECT  0.230 0.000 0.470 1.300 ;
        END
    END VSS
END nd03d2

MACRO nd03d1
    CLASS CORE ;
    FOREIGN nd03d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.390 2.180 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 1.900 ;
        RECT  1.180 1.460 1.490 2.620 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.453  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.220 0.800 2.540 ;
        RECT  0.120 2.220 0.500 3.020 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.885  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.150 3.260 2.680 3.500 ;
        RECT  2.420 1.460 2.680 3.500 ;
        RECT  2.300 1.460 2.680 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  2.190 4.710 2.590 5.600 ;
        RECT  0.870 4.270 1.110 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  0.270 0.000 0.670 0.890 ;
        END
    END VSS
END nd03d1

MACRO nd03d0
    CLASS CORE ;
    FOREIGN nd03d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.100 0.810 2.340 ;
        RECT  0.120 2.100 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 1.900 ;
        RECT  1.180 1.460 1.420 2.380 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.180 3.020 ;
        RECT  1.900 1.980 2.180 3.020 ;
        END
    END A3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.864  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.260 2.680 4.140 ;
        RECT  2.430 1.500 2.680 4.140 ;
        RECT  2.080 1.500 2.680 1.740 ;
        RECT  1.450 3.260 2.680 3.500 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  2.180 4.710 2.580 5.600 ;
        RECT  1.460 4.350 1.700 5.600 ;
        RECT  0.690 3.200 0.930 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  0.160 0.000 0.570 0.890 ;
        END
    END VSS
END nd03d0

MACRO nd02da
    CLASS CORE ;
    FOREIGN nd02da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.462  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.590 3.100 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.180 3.580 ;
        RECT  1.310 2.860 1.980 3.180 ;
        RECT  1.310 2.780 1.710 3.180 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.164  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.580 2.580 8.610 3.450 ;
        RECT  8.180 1.180 8.610 3.450 ;
        RECT  4.730 1.220 8.610 3.450 ;
        RECT  6.700 1.180 7.100 3.450 ;
        RECT  5.220 1.180 5.620 3.450 ;
        RECT  3.740 1.220 8.610 1.720 ;
        RECT  3.740 1.180 4.140 1.720 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  8.220 3.920 8.620 5.600 ;
        RECT  6.920 3.920 7.320 5.600 ;
        RECT  5.620 3.920 6.020 5.600 ;
        RECT  4.320 3.920 4.720 5.600 ;
        RECT  3.020 4.020 3.420 5.600 ;
        RECT  1.500 4.020 1.900 5.600 ;
        RECT  0.150 4.530 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.440 0.000 7.840 0.980 ;
        RECT  5.960 0.000 6.360 0.980 ;
        RECT  4.480 0.000 4.880 0.980 ;
        RECT  3.000 0.000 3.400 1.560 ;
        RECT  1.500 0.000 1.900 1.600 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.490 1.080 1.730 ;
        RECT  0.150 1.410 0.550 1.810 ;
        RECT  0.830 1.490 1.080 2.440 ;
        RECT  0.830 2.200 2.340 2.440 ;
        RECT  1.940 2.150 2.340 2.550 ;
        RECT  0.830 1.490 1.070 4.110 ;
        RECT  0.720 3.710 1.120 4.110 ;
        RECT  2.240 1.180 2.760 1.580 ;
        RECT  2.520 1.750 2.850 1.990 ;
        RECT  2.520 1.180 2.760 1.990 ;
        RECT  2.570 1.950 4.500 2.350 ;
        RECT  2.570 1.950 2.970 3.460 ;
        RECT  2.410 3.120 2.790 4.220 ;
        RECT  2.240 3.820 2.790 4.220 ;
    END
END nd02da

MACRO nd02d7
    CLASS CORE ;
    FOREIGN nd02d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.460  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.590 3.100 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.452  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.180 3.020 ;
        RECT  1.310 2.290 1.980 2.620 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.976  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.390 3.050 7.160 3.450 ;
        RECT  6.660 1.600 7.160 3.450 ;
        RECT  6.660 1.200 7.130 3.450 ;
        RECT  3.770 1.260 7.130 1.500 ;
        RECT  5.250 1.180 5.650 1.580 ;
        RECT  3.770 1.170 4.170 1.590 ;
        RECT  3.390 2.760 3.790 3.450 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.730 3.920 7.130 5.600 ;
        RECT  5.430 3.920 5.830 5.600 ;
        RECT  4.130 3.920 4.530 5.600 ;
        RECT  2.830 3.650 3.230 5.600 ;
        RECT  1.460 4.200 1.860 5.600 ;
        RECT  0.150 4.530 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  5.990 0.000 6.390 0.980 ;
        RECT  4.510 0.000 4.910 0.980 ;
        RECT  3.030 0.000 3.430 0.980 ;
        RECT  1.500 0.000 1.900 1.570 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.490 1.080 1.730 ;
        RECT  0.830 1.490 1.080 2.050 ;
        RECT  0.150 1.400 0.550 1.820 ;
        RECT  0.830 1.810 2.410 2.050 ;
        RECT  0.830 1.490 1.070 4.110 ;
        RECT  0.720 3.710 1.120 4.110 ;
        RECT  2.260 1.170 2.670 1.570 ;
        RECT  2.650 2.110 6.300 2.520 ;
        RECT  2.650 1.280 2.890 3.010 ;
        RECT  2.420 2.770 2.660 3.480 ;
        RECT  2.280 3.240 2.520 4.600 ;
        RECT  2.240 3.910 2.520 4.600 ;
        RECT  2.150 4.200 2.570 4.600 ;
    END
END nd02d7

MACRO nd02d4
    CLASS CORE ;
    FOREIGN nd02d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.580 1.620 3.020 ;
        RECT  1.180 1.680 1.440 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.274  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.600 0.840 2.840 ;
        RECT  0.120 2.020 0.500 2.840 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.750 3.130 5.450 3.370 ;
        RECT  3.680 1.850 5.450 2.090 ;
        RECT  4.530 1.850 4.990 3.370 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.360 4.710 4.770 5.600 ;
        RECT  3.010 4.710 3.410 5.600 ;
        RECT  1.710 4.700 2.110 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.450 0.000 4.690 1.330 ;
        RECT  3.030 0.000 3.270 1.330 ;
        RECT  0.230 0.000 0.470 1.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.450 1.170 2.100 1.410 ;
        RECT  1.860 2.450 2.940 2.690 ;
        RECT  1.860 1.170 2.100 3.500 ;
        RECT  0.920 3.260 2.100 3.500 ;
        RECT  2.410 1.600 3.420 1.840 ;
        RECT  2.410 1.600 2.650 2.160 ;
        RECT  3.180 2.380 3.780 2.620 ;
        RECT  2.410 3.050 2.650 3.640 ;
        RECT  3.180 1.600 3.420 3.640 ;
        RECT  2.410 3.400 3.420 3.640 ;
    END
END nd02d4

MACRO nd02d2
    CLASS CORE ;
    FOREIGN nd02d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.823  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.100 2.020 1.620 2.460 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.600 0.820 2.840 ;
        RECT  0.120 2.020 0.500 2.840 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.852  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.090 2.020 2.740 2.460 ;
        RECT  2.090 3.130 2.600 3.450 ;
        RECT  2.090 1.120 2.330 3.450 ;
        RECT  0.750 3.130 2.600 3.370 ;
        RECT  1.350 1.120 2.330 1.360 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.810 4.700 3.210 5.600 ;
        RECT  1.710 4.290 1.950 5.600 ;
        RECT  0.150 4.700 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.630 0.000 2.870 1.440 ;
        RECT  0.230 0.000 0.470 1.440 ;
        END
    END VSS
END nd02d2

MACRO nd02d1
    CLASS CORE ;
    FOREIGN nd02d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.320 1.620 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.600 0.830 2.840 ;
        RECT  0.120 2.600 0.500 3.580 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.152  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.920 3.260 2.120 3.500 ;
        RECT  1.880 1.460 2.120 3.500 ;
        RECT  1.380 1.830 2.120 2.070 ;
        RECT  1.740 1.460 2.120 2.070 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.240 5.600 ;
        RECT  1.690 4.710 2.090 5.600 ;
        RECT  0.230 4.360 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.240 0.740 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
END nd02d1

MACRO nd02d0
    CLASS CORE ;
    FOREIGN nd02d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.320 1.620 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.600 0.830 2.840 ;
        RECT  0.120 2.600 0.500 3.580 ;
        END
    END A2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.762  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.920 3.260 2.120 3.500 ;
        RECT  1.880 1.460 2.120 3.500 ;
        RECT  1.380 1.830 2.120 2.070 ;
        RECT  1.740 1.460 2.120 2.070 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.240 5.600 ;
        RECT  1.690 4.710 2.090 5.600 ;
        RECT  0.230 4.360 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.240 0.740 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
END nd02d0

MACRO mx08d4
    CLASS CORE ;
    FOREIGN mx08d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.020 2.080 11.250 2.320 ;
        RECT  11.010 1.550 11.250 2.320 ;
        RECT  9.580 2.720 10.650 2.960 ;
        RECT  10.020 2.080 10.260 2.960 ;
        RECT  9.580 2.580 10.020 3.020 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 1.600 10.650 1.840 ;
        RECT  9.020 1.460 9.460 1.900 ;
        END
    END I1
    PIN I2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.470 2.580 8.910 3.020 ;
        RECT  8.410 1.520 8.650 2.970 ;
        RECT  7.670 2.730 8.910 2.970 ;
        END
    END I2
    PIN I3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 1.890 8.070 2.460 ;
        END
    END I3
    PIN I4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.820 6.080 3.140 ;
        RECT  5.840 1.660 6.080 3.140 ;
        RECT  5.580 1.460 5.980 1.860 ;
        RECT  5.100 2.820 5.540 3.580 ;
        END
    END I4
    PIN I5
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.140 5.600 2.540 ;
        RECT  4.540 2.020 5.140 2.540 ;
        END
    END I5
    PIN I6
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.090 1.460 3.330 3.110 ;
        RECT  2.860 2.710 3.300 3.580 ;
        END
    END I6
    PIN I7
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.550 1.760 2.790 2.430 ;
        RECT  2.300 1.460 2.740 2.000 ;
        END
    END I7
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.393  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.290 0.790 2.690 ;
        RECT  0.120 2.290 0.500 3.080 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.275  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.240 2.350 16.740 3.020 ;
        END
    END S1
    PIN S2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.368  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.620 2.820 15.510 3.060 ;
        RECT  14.620 2.580 15.060 3.060 ;
        END
    END S2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.911  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  20.810 1.170 21.050 3.530 ;
        RECT  19.360 2.580 21.050 3.020 ;
        RECT  19.360 1.170 19.760 4.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 21.280 5.600 ;
        RECT  19.970 4.440 20.370 5.600 ;
        RECT  18.490 4.710 18.890 5.600 ;
        RECT  16.450 4.710 16.850 5.600 ;
        RECT  12.000 4.710 12.400 5.600 ;
        RECT  9.290 4.710 9.690 5.600 ;
        RECT  6.700 4.710 7.100 5.600 ;
        RECT  4.240 4.710 4.640 5.600 ;
        RECT  1.990 4.060 2.390 5.600 ;
        RECT  0.720 4.010 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 21.280 0.740 ;
        RECT  19.960 0.000 20.360 0.890 ;
        RECT  18.050 0.000 18.990 0.890 ;
        RECT  15.450 0.000 15.850 1.270 ;
        RECT  11.890 0.000 12.290 0.890 ;
        RECT  9.290 0.000 9.690 0.890 ;
        RECT  6.710 0.000 7.110 0.890 ;
        RECT  4.050 0.000 4.290 1.330 ;
        RECT  1.540 0.000 1.940 1.300 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.270 1.820 ;
        RECT  1.030 2.320 1.480 2.720 ;
        RECT  1.030 1.580 1.270 3.180 ;
        RECT  0.740 2.940 1.270 3.180 ;
        RECT  0.740 2.940 0.980 3.560 ;
        RECT  0.150 3.320 0.980 3.560 ;
        RECT  1.510 1.660 1.960 2.060 ;
        RECT  1.720 2.320 2.190 2.730 ;
        RECT  1.720 1.660 1.960 3.740 ;
        RECT  1.460 3.340 1.960 3.740 ;
        RECT  10.540 1.070 11.730 1.310 ;
        RECT  12.630 1.090 13.050 1.370 ;
        RECT  11.490 1.130 13.050 1.370 ;
        RECT  11.490 1.070 11.730 2.940 ;
        RECT  10.890 2.700 11.730 2.940 ;
        RECT  5.260 0.980 6.470 1.220 ;
        RECT  6.230 1.130 6.560 1.350 ;
        RECT  6.320 1.130 6.560 3.980 ;
        RECT  12.450 3.610 13.680 3.850 ;
        RECT  5.780 3.740 12.690 3.980 ;
        RECT  5.470 3.900 6.010 4.140 ;
        RECT  7.540 1.040 8.340 1.280 ;
        RECT  13.340 1.060 14.920 1.300 ;
        RECT  6.860 1.130 7.790 1.370 ;
        RECT  13.340 1.060 13.580 1.850 ;
        RECT  11.970 1.610 13.580 1.850 ;
        RECT  6.860 1.130 7.100 3.500 ;
        RECT  11.970 1.610 12.210 3.500 ;
        RECT  6.860 3.260 12.210 3.500 ;
        RECT  2.740 0.980 3.810 1.220 ;
        RECT  3.570 0.980 3.810 4.110 ;
        RECT  3.570 3.820 5.150 4.080 ;
        RECT  3.190 3.870 4.140 4.110 ;
        RECT  14.720 3.530 14.960 4.460 ;
        RECT  4.910 3.820 5.150 4.620 ;
        RECT  6.240 4.220 14.970 4.460 ;
        RECT  4.910 4.380 6.470 4.620 ;
        RECT  14.630 2.020 16.000 2.260 ;
        RECT  15.760 2.020 16.000 3.570 ;
        RECT  15.760 3.330 16.330 3.570 ;
        RECT  16.570 1.870 17.430 2.110 ;
        RECT  17.190 1.870 17.430 4.270 ;
        RECT  17.190 3.950 17.630 4.270 ;
        RECT  16.090 0.980 17.820 1.250 ;
        RECT  17.420 1.100 17.910 1.380 ;
        RECT  16.090 0.980 16.330 1.780 ;
        RECT  13.820 1.540 16.330 1.780 ;
        RECT  13.820 1.540 14.060 2.350 ;
        RECT  13.110 2.110 14.060 2.350 ;
        RECT  17.670 1.100 17.910 3.380 ;
        RECT  17.670 3.140 18.330 3.380 ;
        RECT  18.150 1.280 18.390 2.900 ;
        RECT  18.150 2.500 18.820 2.900 ;
        RECT  18.580 2.500 18.820 4.190 ;
        RECT  17.930 3.950 18.820 4.190 ;
    END
END mx08d4

MACRO mx08d2
    CLASS CORE ;
    FOREIGN mx08d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.020 2.080 11.250 2.320 ;
        RECT  11.010 1.550 11.250 2.320 ;
        RECT  9.580 2.720 10.650 2.960 ;
        RECT  10.020 2.080 10.260 2.960 ;
        RECT  9.580 2.580 10.020 3.020 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 1.600 10.650 1.840 ;
        RECT  9.020 1.460 9.460 1.900 ;
        END
    END I1
    PIN I2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.470 2.580 8.910 3.020 ;
        RECT  8.410 1.520 8.650 2.970 ;
        RECT  7.670 2.730 8.910 2.970 ;
        END
    END I2
    PIN I3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 1.890 8.070 2.460 ;
        END
    END I3
    PIN I4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.820 6.080 3.140 ;
        RECT  5.840 1.660 6.080 3.140 ;
        RECT  5.580 1.460 5.980 1.860 ;
        RECT  5.100 2.820 5.540 3.580 ;
        END
    END I4
    PIN I5
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.140 5.600 2.540 ;
        RECT  4.540 2.020 5.140 2.540 ;
        END
    END I5
    PIN I6
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.090 1.460 3.330 3.110 ;
        RECT  2.860 2.710 3.300 3.580 ;
        END
    END I6
    PIN I7
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.550 1.760 2.790 2.430 ;
        RECT  2.300 1.460 2.740 2.000 ;
        END
    END I7
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.393  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.290 0.790 2.690 ;
        RECT  0.120 2.290 0.500 3.080 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.275  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.240 2.340 16.740 3.020 ;
        END
    END S1
    PIN S2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.368  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.620 2.820 15.510 3.060 ;
        RECT  14.620 2.580 15.060 3.060 ;
        END
    END S2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.303  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.580 2.580 20.040 3.020 ;
        RECT  19.580 1.480 20.000 4.100 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.720 5.600 ;
        RECT  20.170 4.440 20.570 5.600 ;
        RECT  18.810 4.710 19.210 5.600 ;
        RECT  16.450 4.710 16.850 5.600 ;
        RECT  12.000 4.710 12.400 5.600 ;
        RECT  9.290 4.710 9.690 5.600 ;
        RECT  6.700 4.710 7.100 5.600 ;
        RECT  4.240 4.710 4.640 5.600 ;
        RECT  1.990 4.060 2.390 5.600 ;
        RECT  0.720 4.010 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.720 0.740 ;
        RECT  20.170 0.000 20.570 0.890 ;
        RECT  18.260 0.000 19.200 0.890 ;
        RECT  15.450 0.000 15.850 1.270 ;
        RECT  11.890 0.000 12.290 0.890 ;
        RECT  9.290 0.000 9.690 0.890 ;
        RECT  6.710 0.000 7.110 0.890 ;
        RECT  4.050 0.000 4.290 1.330 ;
        RECT  1.540 0.000 1.940 1.300 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.270 1.820 ;
        RECT  1.030 2.320 1.480 2.720 ;
        RECT  1.030 1.580 1.270 3.180 ;
        RECT  0.740 2.940 1.270 3.180 ;
        RECT  0.740 2.940 0.980 3.560 ;
        RECT  0.150 3.320 0.980 3.560 ;
        RECT  1.510 1.660 1.960 2.060 ;
        RECT  1.720 2.320 2.190 2.730 ;
        RECT  1.720 1.660 1.960 3.740 ;
        RECT  1.460 3.340 1.960 3.740 ;
        RECT  10.540 1.070 11.730 1.310 ;
        RECT  12.630 1.090 13.050 1.370 ;
        RECT  11.490 1.130 13.050 1.370 ;
        RECT  11.490 1.070 11.730 2.940 ;
        RECT  10.890 2.700 11.730 2.940 ;
        RECT  5.260 0.980 6.470 1.220 ;
        RECT  6.230 1.130 6.560 1.350 ;
        RECT  6.320 1.130 6.560 3.980 ;
        RECT  12.450 3.610 13.680 3.850 ;
        RECT  5.780 3.740 12.690 3.980 ;
        RECT  5.470 3.900 6.010 4.140 ;
        RECT  7.540 1.040 8.340 1.280 ;
        RECT  13.340 1.060 14.920 1.300 ;
        RECT  6.860 1.130 7.790 1.370 ;
        RECT  13.340 1.060 13.580 1.850 ;
        RECT  11.970 1.610 13.580 1.850 ;
        RECT  6.860 1.130 7.100 3.500 ;
        RECT  11.970 1.610 12.210 3.500 ;
        RECT  6.860 3.260 12.210 3.500 ;
        RECT  2.740 0.980 3.810 1.220 ;
        RECT  3.570 0.980 3.810 4.110 ;
        RECT  3.570 3.820 5.150 4.080 ;
        RECT  3.190 3.870 4.140 4.110 ;
        RECT  14.720 3.530 14.960 4.460 ;
        RECT  4.910 3.820 5.150 4.620 ;
        RECT  6.240 4.220 14.970 4.460 ;
        RECT  4.910 4.380 6.470 4.620 ;
        RECT  14.630 2.020 16.000 2.260 ;
        RECT  15.760 2.020 16.000 3.570 ;
        RECT  15.760 3.330 16.330 3.570 ;
        RECT  17.240 1.740 17.560 2.060 ;
        RECT  16.570 1.820 17.560 2.060 ;
        RECT  17.240 1.740 17.480 3.650 ;
        RECT  17.230 3.250 17.630 3.650 ;
        RECT  16.090 0.980 17.980 1.250 ;
        RECT  17.520 1.150 18.050 1.440 ;
        RECT  16.090 0.980 16.330 1.780 ;
        RECT  13.820 1.540 16.330 1.780 ;
        RECT  13.820 1.540 14.060 2.400 ;
        RECT  13.190 2.160 14.060 2.400 ;
        RECT  17.810 2.710 18.240 2.950 ;
        RECT  17.810 1.150 18.050 2.950 ;
        RECT  18.010 2.720 18.250 3.460 ;
        RECT  18.290 1.610 18.740 2.010 ;
        RECT  18.500 1.610 18.740 4.430 ;
        RECT  17.930 4.190 18.740 4.430 ;
    END
END mx08d2

MACRO mx08d1
    CLASS CORE ;
    FOREIGN mx08d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.020 2.080 11.250 2.320 ;
        RECT  11.010 1.550 11.250 2.320 ;
        RECT  9.580 2.720 10.650 2.960 ;
        RECT  10.020 2.080 10.260 2.960 ;
        RECT  9.580 2.580 10.020 3.020 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 1.600 10.650 1.840 ;
        RECT  9.020 1.460 9.460 1.900 ;
        END
    END I1
    PIN I2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.470 2.580 8.910 3.020 ;
        RECT  8.410 1.520 8.650 2.970 ;
        RECT  7.670 2.730 8.910 2.970 ;
        END
    END I2
    PIN I3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 1.890 8.070 2.460 ;
        END
    END I3
    PIN I4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.900 6.080 3.140 ;
        RECT  5.840 1.660 6.080 3.140 ;
        RECT  5.580 1.460 5.980 1.860 ;
        RECT  5.100 2.900 5.540 3.580 ;
        RECT  5.100 2.820 5.530 3.580 ;
        END
    END I4
    PIN I5
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.140 5.600 2.540 ;
        RECT  4.540 2.020 5.140 2.540 ;
        END
    END I5
    PIN I6
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.090 1.460 3.330 3.110 ;
        RECT  2.850 2.710 3.300 3.580 ;
        END
    END I6
    PIN I7
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.550 1.760 2.790 2.430 ;
        RECT  2.300 1.460 2.740 2.000 ;
        END
    END I7
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.393  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.290 0.790 2.690 ;
        RECT  0.120 2.290 0.500 3.080 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.275  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.240 2.340 16.740 3.020 ;
        END
    END S1
    PIN S2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.368  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.620 2.820 15.510 3.060 ;
        RECT  14.620 2.580 15.060 3.060 ;
        END
    END S2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.250  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.600 2.580 20.040 3.020 ;
        RECT  19.600 1.480 20.000 4.560 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.160 5.600 ;
        RECT  18.810 4.710 19.210 5.600 ;
        RECT  16.450 4.710 16.850 5.600 ;
        RECT  12.000 4.710 12.400 5.600 ;
        RECT  9.290 4.710 9.690 5.600 ;
        RECT  6.700 4.710 7.100 5.600 ;
        RECT  4.240 4.710 4.640 5.600 ;
        RECT  1.990 4.060 2.390 5.600 ;
        RECT  0.720 4.010 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.160 0.740 ;
        RECT  18.290 0.000 19.230 1.200 ;
        RECT  15.450 0.000 15.850 1.270 ;
        RECT  11.890 0.000 12.290 0.890 ;
        RECT  9.290 0.000 9.690 0.890 ;
        RECT  6.710 0.000 7.110 0.890 ;
        RECT  4.050 0.000 4.290 1.330 ;
        RECT  1.540 0.000 1.940 1.300 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.270 1.820 ;
        RECT  1.030 2.320 1.480 2.720 ;
        RECT  1.030 1.580 1.270 3.180 ;
        RECT  0.740 2.940 1.270 3.180 ;
        RECT  0.740 2.940 0.980 3.560 ;
        RECT  0.150 3.320 0.980 3.560 ;
        RECT  1.510 1.660 1.960 2.060 ;
        RECT  1.720 2.320 2.190 2.730 ;
        RECT  1.720 1.660 1.960 3.740 ;
        RECT  1.460 3.340 1.960 3.740 ;
        RECT  10.540 1.070 11.730 1.310 ;
        RECT  12.630 1.090 13.050 1.370 ;
        RECT  11.490 1.130 13.050 1.370 ;
        RECT  11.490 1.070 11.730 2.940 ;
        RECT  10.890 2.700 11.730 2.940 ;
        RECT  5.260 0.980 6.470 1.220 ;
        RECT  6.230 1.130 6.560 1.350 ;
        RECT  6.320 1.130 6.560 3.980 ;
        RECT  12.450 3.610 13.680 3.850 ;
        RECT  5.800 3.740 12.690 3.980 ;
        RECT  5.470 3.860 6.010 4.100 ;
        RECT  7.540 1.040 8.340 1.280 ;
        RECT  13.340 1.060 14.920 1.300 ;
        RECT  6.860 1.130 7.790 1.370 ;
        RECT  13.340 1.060 13.580 1.850 ;
        RECT  11.970 1.610 13.580 1.850 ;
        RECT  6.860 1.130 7.100 3.500 ;
        RECT  11.970 1.610 12.210 3.500 ;
        RECT  6.860 3.260 12.210 3.500 ;
        RECT  2.740 0.980 3.810 1.220 ;
        RECT  3.570 0.980 3.810 4.110 ;
        RECT  3.570 3.820 5.150 4.080 ;
        RECT  3.190 3.870 4.140 4.110 ;
        RECT  14.720 3.530 14.960 4.460 ;
        RECT  4.910 3.820 5.150 4.620 ;
        RECT  6.240 4.220 14.970 4.460 ;
        RECT  4.910 4.380 6.470 4.620 ;
        RECT  14.630 2.020 16.000 2.260 ;
        RECT  15.760 2.020 16.000 3.570 ;
        RECT  15.760 3.330 16.330 3.570 ;
        RECT  17.240 1.740 17.560 2.060 ;
        RECT  16.570 1.820 17.560 2.060 ;
        RECT  17.240 1.740 17.480 3.650 ;
        RECT  17.230 3.250 17.630 3.650 ;
        RECT  16.090 0.980 18.050 1.250 ;
        RECT  17.520 0.980 18.050 1.440 ;
        RECT  16.090 0.980 16.330 1.780 ;
        RECT  13.820 1.540 16.330 1.780 ;
        RECT  13.820 1.540 14.060 2.330 ;
        RECT  13.110 2.090 14.060 2.330 ;
        RECT  17.810 2.710 18.240 2.950 ;
        RECT  17.810 0.980 18.050 2.950 ;
        RECT  18.010 2.720 18.250 3.460 ;
        RECT  18.310 1.610 18.740 2.010 ;
        RECT  18.500 1.610 18.740 4.430 ;
        RECT  17.930 4.190 18.740 4.430 ;
    END
END mx08d1

MACRO mx04d4
    CLASS CORE ;
    FOREIGN mx04d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.690 2.530 3.300 3.020 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.300 2.250 6.580 3.020 ;
        RECT  6.070 2.250 6.580 2.650 ;
        END
    END I1
    PIN I2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.180 6.100 3.510 ;
        END
    END I2
    PIN I3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.650 2.580 9.460 3.020 ;
        END
    END I3
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.035  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.630 3.850 7.830 4.090 ;
        RECT  7.590 1.920 7.830 4.090 ;
        RECT  4.060 3.750 6.870 3.990 ;
        RECT  1.510 3.850 4.420 4.090 ;
        RECT  4.060 3.140 4.420 4.090 ;
        RECT  1.510 3.210 1.970 4.090 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.581  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.450 2.100 5.540 2.410 ;
        RECT  3.540 2.650 4.690 2.890 ;
        RECT  4.450 2.100 4.690 2.890 ;
        RECT  2.210 3.280 3.820 3.610 ;
        RECT  3.540 2.650 3.820 3.610 ;
        RECT  2.210 2.600 2.450 3.610 ;
        RECT  1.190 2.600 2.450 2.880 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.870 3.460 13.590 3.860 ;
        RECT  11.860 1.720 13.590 2.120 ;
        RECT  12.940 1.720 13.380 3.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 14.000 5.600 ;
        RECT  12.520 4.150 12.760 5.600 ;
        RECT  11.210 4.150 11.450 5.600 ;
        RECT  8.980 4.380 9.220 5.600 ;
        RECT  5.550 4.710 5.950 5.600 ;
        RECT  2.210 4.380 2.550 5.600 ;
        RECT  0.230 4.050 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 14.000 0.740 ;
        RECT  12.680 0.000 12.920 1.420 ;
        RECT  11.380 0.000 11.620 1.420 ;
        RECT  9.190 0.000 9.590 0.890 ;
        RECT  5.810 0.000 6.210 0.890 ;
        RECT  2.430 0.000 2.830 0.990 ;
        RECT  1.220 0.000 1.490 1.880 ;
        RECT  0.470 0.000 0.960 0.830 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.620 0.830 1.860 ;
        RECT  0.230 1.620 0.470 3.460 ;
        RECT  1.860 1.610 7.340 1.850 ;
        RECT  1.860 1.390 2.180 2.360 ;
        RECT  0.710 2.120 2.180 2.360 ;
        RECT  3.950 1.610 4.190 2.410 ;
        RECT  7.100 1.610 7.340 3.610 ;
        RECT  0.710 2.120 0.950 4.620 ;
        RECT  0.710 4.360 1.840 4.620 ;
        RECT  4.120 0.980 5.570 1.220 ;
        RECT  5.300 1.130 8.340 1.370 ;
        RECT  8.100 2.000 9.790 2.240 ;
        RECT  5.110 4.230 6.390 4.470 ;
        RECT  3.850 4.330 5.350 4.570 ;
        RECT  8.100 1.130 8.340 4.570 ;
        RECT  6.150 4.330 8.340 4.570 ;
        RECT  9.760 1.230 10.270 1.640 ;
        RECT  10.030 2.250 11.130 2.650 ;
        RECT  10.030 1.230 10.270 4.520 ;
        RECT  9.580 4.110 10.270 4.520 ;
        RECT  10.560 1.660 11.610 1.900 ;
        RECT  11.370 2.360 12.550 2.760 ;
        RECT  11.370 1.660 11.610 3.200 ;
        RECT  10.630 2.960 11.610 3.200 ;
        RECT  10.630 2.960 10.900 3.590 ;
    END
END mx04d4

MACRO mx04d2
    CLASS CORE ;
    FOREIGN mx04d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.690 2.530 3.300 3.020 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.300 2.310 6.580 3.020 ;
        RECT  6.070 2.310 6.580 2.660 ;
        END
    END I1
    PIN I2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.401  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.270 3.220 6.100 3.500 ;
        END
    END I2
    PIN I3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.650 2.580 9.460 3.020 ;
        END
    END I3
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.057  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.630 3.850 7.830 4.090 ;
        RECT  7.590 1.960 7.830 4.090 ;
        RECT  4.100 3.750 6.870 3.990 ;
        RECT  1.510 3.780 4.420 4.070 ;
        RECT  4.100 3.210 4.420 4.070 ;
        RECT  1.510 3.210 1.970 4.070 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.540 2.650 5.250 2.940 ;
        RECT  4.950 2.090 5.250 2.940 ;
        RECT  2.210 3.280 3.820 3.540 ;
        RECT  3.540 2.650 3.820 3.540 ;
        RECT  2.210 2.600 2.450 3.540 ;
        RECT  1.190 2.600 2.450 2.880 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.273  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.580 3.300 10.270 4.140 ;
        RECT  10.030 1.430 10.270 4.140 ;
        RECT  9.770 1.430 10.270 1.800 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.760 5.600 ;
        RECT  10.330 4.380 10.570 5.600 ;
        RECT  8.980 4.380 9.220 5.600 ;
        RECT  5.550 4.710 5.950 5.600 ;
        RECT  2.210 4.380 2.550 5.600 ;
        RECT  0.230 4.050 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.760 0.740 ;
        RECT  10.580 0.000 10.830 1.210 ;
        RECT  9.190 0.000 9.500 1.210 ;
        RECT  5.810 0.000 6.210 0.890 ;
        RECT  2.430 0.000 2.830 0.990 ;
        RECT  1.220 0.000 1.490 1.880 ;
        RECT  0.470 0.000 0.960 0.830 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.620 0.830 1.860 ;
        RECT  0.230 1.620 0.470 3.460 ;
        RECT  1.860 1.610 7.340 1.850 ;
        RECT  1.860 1.390 2.180 2.360 ;
        RECT  0.710 2.120 2.180 2.360 ;
        RECT  3.950 1.610 4.190 2.410 ;
        RECT  7.100 1.610 7.340 3.610 ;
        RECT  0.710 2.120 0.950 4.620 ;
        RECT  0.710 4.360 1.840 4.620 ;
        RECT  4.120 0.980 5.570 1.220 ;
        RECT  6.480 0.980 8.340 1.290 ;
        RECT  5.300 1.130 6.720 1.370 ;
        RECT  8.100 2.060 9.790 2.310 ;
        RECT  5.110 4.230 6.390 4.470 ;
        RECT  3.850 4.330 5.350 4.570 ;
        RECT  8.100 0.980 8.340 4.570 ;
        RECT  6.150 4.330 8.340 4.570 ;
    END
END mx04d2

MACRO mx04d1
    CLASS CORE ;
    FOREIGN mx04d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.690 2.530 3.300 3.020 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.300 2.250 6.580 3.020 ;
        RECT  6.070 2.250 6.580 2.650 ;
        END
    END I1
    PIN I2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.270 3.220 6.100 3.510 ;
        RECT  5.270 3.100 5.740 3.510 ;
        END
    END I2
    PIN I3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.650 2.580 9.460 3.020 ;
        END
    END I3
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.035  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.630 3.850 7.830 4.090 ;
        RECT  7.590 1.920 7.830 4.090 ;
        RECT  4.060 3.750 6.870 3.990 ;
        RECT  1.510 3.850 4.420 4.090 ;
        RECT  4.060 3.140 4.420 4.090 ;
        RECT  1.510 3.210 1.970 4.090 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.581  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.450 2.100 5.540 2.410 ;
        RECT  3.540 2.650 4.690 2.890 ;
        RECT  4.450 2.100 4.690 2.890 ;
        RECT  2.210 3.280 3.820 3.610 ;
        RECT  3.540 2.650 3.820 3.610 ;
        RECT  2.210 2.600 2.450 3.610 ;
        RECT  1.190 2.600 2.450 2.880 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.163  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.580 3.700 10.270 4.520 ;
        RECT  10.030 1.360 10.270 4.520 ;
        RECT  9.820 1.360 10.270 1.770 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  8.980 4.380 9.220 5.600 ;
        RECT  5.550 4.710 5.950 5.600 ;
        RECT  2.210 4.380 2.550 5.600 ;
        RECT  0.230 4.050 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  9.190 0.000 9.590 0.890 ;
        RECT  5.810 0.000 6.210 0.890 ;
        RECT  2.430 0.000 2.830 0.990 ;
        RECT  1.220 0.000 1.490 1.880 ;
        RECT  0.470 0.000 0.960 0.830 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.620 0.830 1.860 ;
        RECT  0.230 1.620 0.470 3.460 ;
        RECT  1.860 1.610 7.340 1.850 ;
        RECT  1.860 1.390 2.180 2.360 ;
        RECT  0.710 2.120 2.180 2.360 ;
        RECT  3.950 1.610 4.190 2.410 ;
        RECT  7.100 1.610 7.340 3.610 ;
        RECT  0.710 2.120 0.950 4.620 ;
        RECT  0.710 4.360 1.840 4.620 ;
        RECT  4.120 0.980 5.570 1.220 ;
        RECT  5.300 1.130 8.340 1.370 ;
        RECT  8.100 2.010 9.790 2.250 ;
        RECT  5.110 4.230 6.390 4.470 ;
        RECT  3.850 4.330 5.350 4.570 ;
        RECT  8.100 1.130 8.340 4.570 ;
        RECT  6.150 4.330 8.340 4.570 ;
    END
END mx04d1

MACRO mx04d0
    CLASS CORE ;
    FOREIGN mx04d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.690 2.530 3.300 3.020 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.300 2.250 6.580 3.020 ;
        RECT  6.070 2.250 6.580 2.650 ;
        END
    END I1
    PIN I2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.270 3.220 6.100 3.510 ;
        RECT  5.270 3.100 5.740 3.510 ;
        END
    END I2
    PIN I3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.650 2.580 9.460 3.020 ;
        END
    END I3
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.035  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.630 3.850 7.830 4.090 ;
        RECT  7.590 1.920 7.830 4.090 ;
        RECT  4.060 3.750 6.870 3.990 ;
        RECT  1.510 3.850 4.420 4.090 ;
        RECT  4.060 3.140 4.420 4.090 ;
        RECT  1.510 3.210 1.970 4.090 ;
        END
    END S0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.581  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.450 2.100 5.540 2.410 ;
        RECT  3.540 2.650 4.690 2.890 ;
        RECT  4.450 2.100 4.690 2.890 ;
        RECT  2.210 3.280 3.820 3.610 ;
        RECT  3.540 2.650 3.820 3.610 ;
        RECT  2.210 2.600 2.450 3.610 ;
        RECT  1.190 2.600 2.450 2.880 ;
        END
    END S1
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.617  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.580 3.700 10.270 4.520 ;
        RECT  10.030 1.230 10.270 4.520 ;
        RECT  9.760 1.230 10.270 1.640 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  8.980 4.380 9.220 5.600 ;
        RECT  5.550 4.710 5.950 5.600 ;
        RECT  2.210 4.380 2.550 5.600 ;
        RECT  0.230 4.050 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  9.190 0.000 9.590 0.890 ;
        RECT  5.810 0.000 6.210 0.890 ;
        RECT  2.430 0.000 2.830 0.990 ;
        RECT  1.220 0.000 1.490 1.880 ;
        RECT  0.470 0.000 0.960 0.830 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.620 0.830 1.860 ;
        RECT  0.230 1.620 0.470 3.460 ;
        RECT  1.860 1.610 7.340 1.850 ;
        RECT  1.860 1.390 2.180 2.360 ;
        RECT  0.710 2.120 2.180 2.360 ;
        RECT  3.950 1.610 4.190 2.410 ;
        RECT  7.100 1.610 7.340 3.610 ;
        RECT  0.710 2.120 0.950 4.620 ;
        RECT  0.710 4.360 1.840 4.620 ;
        RECT  4.120 0.980 5.570 1.220 ;
        RECT  5.300 1.130 8.340 1.370 ;
        RECT  8.100 2.000 9.790 2.240 ;
        RECT  5.110 4.230 6.390 4.470 ;
        RECT  3.850 4.330 5.350 4.570 ;
        RECT  8.100 1.130 8.340 4.570 ;
        RECT  6.150 4.330 8.340 4.570 ;
    END
END mx04d0

MACRO mx02d4
    CLASS CORE ;
    FOREIGN mx02d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.474  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.820 2.020 3.220 2.650 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.260 1.540 3.020 ;
        END
    END I1
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.170 0.460 3.020 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.329  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.740 3.460 5.460 3.860 ;
        RECT  5.180 1.720 5.460 3.860 ;
        RECT  3.730 1.720 5.460 2.120 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.390 4.150 4.630 5.600 ;
        RECT  3.080 4.150 3.320 5.600 ;
        RECT  0.720 4.180 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.550 0.000 4.790 1.420 ;
        RECT  3.250 0.000 3.490 1.420 ;
        RECT  0.720 0.000 1.120 0.900 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.480 0.940 1.720 ;
        RECT  0.700 1.690 2.100 1.930 ;
        RECT  1.860 1.690 2.100 2.940 ;
        RECT  0.700 1.480 0.940 3.500 ;
        RECT  0.150 3.260 0.940 3.500 ;
        RECT  1.970 1.020 2.580 1.420 ;
        RECT  3.480 2.360 4.420 2.760 ;
        RECT  2.340 2.960 3.800 3.200 ;
        RECT  3.480 2.360 3.800 3.200 ;
        RECT  2.340 1.020 2.580 3.580 ;
        RECT  1.940 3.180 2.580 3.580 ;
    END
END mx02d4

MACRO mx02d2
    CLASS CORE ;
    FOREIGN mx02d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.474  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.820 2.020 3.220 2.650 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.520 1.540 3.160 ;
        END
    END I1
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.170 0.460 3.020 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.195  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.800 3.460 4.420 3.860 ;
        RECT  3.980 3.140 4.420 3.860 ;
        RECT  3.980 1.800 4.220 3.860 ;
        RECT  3.710 1.800 4.220 2.040 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.450 4.150 4.690 5.600 ;
        RECT  3.140 4.150 3.380 5.600 ;
        RECT  0.720 4.180 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.530 0.000 4.770 1.420 ;
        RECT  3.230 0.000 3.470 1.420 ;
        RECT  0.720 0.000 1.120 1.110 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.690 2.100 1.930 ;
        RECT  1.860 1.690 2.100 2.940 ;
        RECT  0.700 1.690 0.940 3.500 ;
        RECT  0.150 3.260 0.940 3.500 ;
        RECT  1.950 1.020 2.580 1.420 ;
        RECT  2.340 2.960 3.740 3.200 ;
        RECT  3.500 2.280 3.740 3.200 ;
        RECT  2.340 1.020 2.580 3.580 ;
        RECT  2.020 3.180 2.580 3.580 ;
    END
END mx02d2

MACRO mx02d1
    CLASS CORE ;
    FOREIGN mx02d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.449  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.910 1.970 3.280 2.570 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.250 2.520 1.580 3.160 ;
        END
    END I1
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.170 0.530 3.020 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.134  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.010 3.520 4.360 4.260 ;
        RECT  4.120 1.720 4.360 4.260 ;
        RECT  3.930 1.720 4.360 1.960 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.270 4.090 3.510 5.600 ;
        RECT  0.970 4.090 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.370 0.000 3.610 1.420 ;
        RECT  0.860 0.000 1.260 1.110 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.650 2.170 1.890 ;
        RECT  1.930 1.650 2.170 2.940 ;
        RECT  0.770 1.650 1.010 3.620 ;
        RECT  0.230 3.380 1.010 3.620 ;
        RECT  0.230 3.380 0.470 4.280 ;
        RECT  2.090 1.100 2.670 1.340 ;
        RECT  3.640 2.220 3.880 3.170 ;
        RECT  2.430 2.930 3.880 3.170 ;
        RECT  2.430 1.100 2.670 3.490 ;
        RECT  2.090 3.250 2.670 3.490 ;
    END
END mx02d1

MACRO mx02d0
    CLASS CORE ;
    FOREIGN mx02d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.281  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 2.580 3.280 3.380 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.580 1.540 3.210 ;
        END
    END I1
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.580 0.460 3.530 ;
        END
    END S
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.887  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.930 4.100 4.340 4.420 ;
        RECT  4.060 1.320 4.340 4.420 ;
        RECT  3.930 1.320 4.340 1.720 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  2.960 4.710 3.360 5.600 ;
        RECT  1.160 4.510 1.560 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.160 0.000 3.560 0.890 ;
        RECT  0.800 0.000 1.200 1.310 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.210 1.710 0.610 2.110 ;
        RECT  0.210 1.870 2.100 2.110 ;
        RECT  1.860 1.870 2.100 3.250 ;
        RECT  0.700 1.870 0.940 4.170 ;
        RECT  0.210 3.770 0.940 4.170 ;
        RECT  2.030 1.390 3.000 1.630 ;
        RECT  2.760 1.390 3.000 2.190 ;
        RECT  2.760 1.950 3.760 2.190 ;
        RECT  3.520 1.950 3.760 3.860 ;
        RECT  2.030 3.620 3.760 3.860 ;
    END
END mx02d0

MACRO mi02d4
    CLASS CORE ;
    FOREIGN mi02d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.920 2.690 3.220 3.580 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.390 1.540 3.580 ;
        END
    END I1
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.050 0.520 3.110 ;
        END
    END S
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.378  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.040 3.050 6.750 3.450 ;
        RECT  6.410 1.620 6.750 3.450 ;
        RECT  5.040 1.620 6.750 2.020 ;
        RECT  5.040 3.050 5.540 4.140 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  5.610 4.540 6.010 5.600 ;
        RECT  4.270 4.540 4.670 5.600 ;
        RECT  3.120 4.710 3.520 5.600 ;
        RECT  0.800 4.160 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  5.610 0.000 6.010 1.330 ;
        RECT  4.300 0.000 4.700 1.330 ;
        RECT  3.200 0.000 3.440 1.330 ;
        RECT  0.720 0.000 1.120 1.200 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.570 2.200 1.810 ;
        RECT  1.960 1.570 2.200 3.010 ;
        RECT  0.760 1.570 1.000 3.790 ;
        RECT  0.150 3.550 1.000 3.790 ;
        RECT  1.920 1.090 2.680 1.330 ;
        RECT  2.440 2.210 3.640 2.450 ;
        RECT  3.460 2.230 3.930 2.630 ;
        RECT  2.440 1.090 2.680 4.440 ;
        RECT  1.920 4.200 2.680 4.440 ;
        RECT  3.750 1.750 4.460 1.990 ;
        RECT  4.220 2.410 5.160 2.810 ;
        RECT  4.220 1.750 4.460 3.790 ;
        RECT  3.770 3.550 4.460 3.790 ;
    END
END mi02d4

MACRO mi02d2
    CLASS CORE ;
    FOREIGN mi02d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.920 2.690 3.220 3.580 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.390 1.540 3.580 ;
        END
    END I1
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.050 0.520 3.110 ;
        END
    END S
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.179  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.120 1.620 5.460 3.450 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.690 4.090 5.930 5.600 ;
        RECT  4.350 4.340 4.590 5.600 ;
        RECT  3.140 4.710 3.540 5.600 ;
        RECT  0.800 4.160 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.610 0.000 6.010 1.330 ;
        RECT  4.300 0.000 4.700 1.330 ;
        RECT  3.200 0.000 3.440 1.330 ;
        RECT  0.720 0.000 1.120 1.200 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.570 2.200 1.810 ;
        RECT  1.960 1.570 2.200 3.010 ;
        RECT  0.760 1.570 1.000 3.790 ;
        RECT  0.150 3.550 1.000 3.790 ;
        RECT  1.920 1.090 2.680 1.330 ;
        RECT  2.440 2.210 3.640 2.450 ;
        RECT  3.460 2.230 3.930 2.630 ;
        RECT  2.440 1.090 2.680 4.440 ;
        RECT  1.920 4.200 2.680 4.440 ;
        RECT  3.750 1.750 4.460 1.990 ;
        RECT  4.220 2.210 4.620 2.610 ;
        RECT  4.220 1.750 4.460 3.790 ;
        RECT  3.770 3.550 4.460 3.790 ;
    END
END mi02d2

MACRO mi02d1
    CLASS CORE ;
    FOREIGN mi02d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.920 2.700 3.220 3.580 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.390 1.540 3.580 ;
        END
    END I1
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.050 0.520 3.110 ;
        END
    END S
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.019  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.130 1.620 5.460 4.140 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.560 4.130 4.800 5.600 ;
        RECT  3.000 4.580 3.400 5.600 ;
        RECT  0.800 4.160 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.480 0.000 4.880 1.330 ;
        RECT  3.200 0.000 3.440 1.330 ;
        RECT  0.720 0.000 1.120 1.200 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.570 2.200 1.810 ;
        RECT  1.960 1.570 2.200 3.010 ;
        RECT  0.760 1.570 1.000 3.790 ;
        RECT  0.150 3.550 1.000 3.790 ;
        RECT  1.920 1.090 2.680 1.330 ;
        RECT  2.440 2.220 3.620 2.460 ;
        RECT  3.450 2.230 3.930 2.630 ;
        RECT  2.440 1.090 2.680 4.440 ;
        RECT  1.920 4.200 2.680 4.440 ;
        RECT  3.750 1.750 4.460 1.990 ;
        RECT  4.220 2.210 4.620 2.610 ;
        RECT  4.220 1.750 4.460 3.790 ;
        RECT  3.780 3.550 4.460 3.790 ;
    END
END mi02d1

MACRO mi02d0
    CLASS CORE ;
    FOREIGN mi02d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.900 3.140 3.440 3.580 ;
        RECT  3.200 2.710 3.440 3.580 ;
        END
    END I0
    PIN I1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 3.140 2.180 3.580 ;
        RECT  1.260 2.710 1.660 3.580 ;
        END
    END I1
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.050 0.540 3.110 ;
        END
    END S
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.835  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.130 1.550 5.460 4.620 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.270 4.620 4.670 5.600 ;
        RECT  3.090 4.350 3.490 5.600 ;
        RECT  0.820 4.160 1.060 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  3.320 0.000 3.560 1.870 ;
        RECT  0.820 0.000 1.060 1.030 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.570 2.480 1.810 ;
        RECT  2.240 1.570 2.480 2.420 ;
        RECT  0.780 1.570 1.020 3.590 ;
        RECT  0.170 3.350 1.020 3.590 ;
        RECT  1.970 1.090 2.960 1.330 ;
        RECT  2.720 2.110 3.830 2.350 ;
        RECT  2.720 1.090 2.960 2.900 ;
        RECT  2.420 2.660 2.960 2.900 ;
        RECT  2.420 2.660 2.660 4.190 ;
        RECT  2.010 3.950 2.660 4.190 ;
        RECT  3.980 1.490 4.380 1.890 ;
        RECT  4.140 2.030 4.640 2.430 ;
        RECT  4.140 1.490 4.380 3.640 ;
        RECT  4.050 3.240 4.450 3.640 ;
    END
END mi02d0

MACRO mffnrb4
    CLASS CORE ;
    FOREIGN mffnrb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.600 2.480 6.190 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.384  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 1.910 2.780 2.460 ;
        RECT  2.270 1.910 2.590 2.880 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.380  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.380 0.980 2.620 ;
        RECT  0.130 2.380 0.500 3.030 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.257  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  20.780 1.370 21.510 1.900 ;
        RECT  18.940 3.370 21.120 3.770 ;
        RECT  20.780 1.370 21.120 3.770 ;
        RECT  19.570 1.370 21.510 1.770 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.187  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.730 1.450 18.700 1.690 ;
        RECT  17.440 1.450 17.900 1.900 ;
        RECT  17.440 2.970 17.870 3.370 ;
        RECT  16.080 3.630 17.680 3.870 ;
        RECT  17.440 1.450 17.680 3.870 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 21.840 5.600 ;
        RECT  21.050 4.320 21.450 5.600 ;
        RECT  19.710 4.320 20.110 5.600 ;
        RECT  18.410 4.180 18.650 5.600 ;
        RECT  16.770 4.590 17.170 5.600 ;
        RECT  15.380 4.590 15.780 5.600 ;
        RECT  14.580 4.680 14.980 5.600 ;
        RECT  13.080 4.340 13.480 5.600 ;
        RECT  9.830 4.710 10.230 5.600 ;
        RECT  6.410 4.710 6.830 5.600 ;
        RECT  5.000 4.710 5.400 5.600 ;
        RECT  2.230 4.220 2.610 5.600 ;
        RECT  0.760 4.330 1.160 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 21.840 0.740 ;
        RECT  20.340 0.000 20.740 1.130 ;
        RECT  18.800 0.000 19.200 0.890 ;
        RECT  17.500 0.000 17.900 0.900 ;
        RECT  15.960 0.000 16.360 0.890 ;
        RECT  13.680 0.000 14.080 0.890 ;
        RECT  10.940 0.000 11.180 1.850 ;
        RECT  7.080 0.000 7.480 0.890 ;
        RECT  5.630 0.000 5.870 1.840 ;
        RECT  1.990 0.000 2.390 0.890 ;
        RECT  1.020 0.000 1.420 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 0.980 0.460 2.090 ;
        RECT  0.180 1.290 0.590 2.090 ;
        RECT  0.180 1.850 1.460 2.090 ;
        RECT  1.220 1.850 1.460 3.510 ;
        RECT  0.260 3.270 1.460 3.510 ;
        RECT  0.260 3.270 0.500 3.930 ;
        RECT  3.040 1.560 3.280 2.360 ;
        RECT  3.020 2.120 3.260 3.500 ;
        RECT  2.760 3.100 3.260 3.500 ;
        RECT  2.620 0.980 4.500 1.220 ;
        RECT  1.770 1.160 2.860 1.400 ;
        RECT  1.770 1.160 2.010 3.410 ;
        RECT  1.820 3.170 2.060 3.980 ;
        RECT  1.820 3.740 3.740 3.980 ;
        RECT  3.500 2.520 3.740 3.980 ;
        RECT  1.500 3.790 2.010 4.030 ;
        RECT  4.460 1.590 5.200 1.830 ;
        RECT  4.460 1.590 4.700 3.510 ;
        RECT  6.110 0.980 6.490 1.960 ;
        RECT  6.110 1.390 6.570 1.960 ;
        RECT  6.110 1.510 6.900 1.960 ;
        RECT  6.660 1.510 6.900 3.500 ;
        RECT  5.730 3.260 6.900 3.500 ;
        RECT  5.730 3.260 5.970 3.820 ;
        RECT  8.380 1.550 8.930 1.790 ;
        RECT  8.380 1.550 8.620 2.280 ;
        RECT  7.930 2.040 8.620 2.280 ;
        RECT  3.980 1.540 4.220 4.460 ;
        RECT  3.590 4.220 4.970 4.460 ;
        RECT  3.980 4.160 4.970 4.460 ;
        RECT  7.930 2.040 8.170 4.470 ;
        RECT  4.540 4.230 8.170 4.470 ;
        RECT  7.800 0.980 10.000 1.220 ;
        RECT  7.800 0.980 8.040 1.790 ;
        RECT  7.380 1.550 8.040 1.790 ;
        RECT  7.380 1.550 7.620 3.980 ;
        RECT  6.980 3.740 7.620 3.980 ;
        RECT  9.990 1.460 10.490 1.860 ;
        RECT  9.990 1.460 10.230 2.280 ;
        RECT  9.650 2.040 10.230 2.280 ;
        RECT  9.650 2.040 9.890 3.990 ;
        RECT  9.330 3.750 9.890 3.990 ;
        RECT  9.170 1.560 9.750 1.800 ;
        RECT  9.170 1.560 9.410 2.380 ;
        RECT  9.010 2.140 9.250 2.760 ;
        RECT  8.670 2.520 9.250 2.760 ;
        RECT  8.670 2.520 8.910 4.470 ;
        RECT  10.660 3.100 10.900 4.470 ;
        RECT  8.670 4.230 10.900 4.470 ;
        RECT  11.680 1.470 11.920 2.350 ;
        RECT  10.470 2.110 11.920 2.350 ;
        RECT  11.200 2.110 11.440 3.550 ;
        RECT  13.580 1.130 15.930 1.370 ;
        RECT  15.690 1.130 15.930 1.690 ;
        RECT  13.580 1.130 13.820 1.760 ;
        RECT  12.910 1.520 13.820 1.760 ;
        RECT  12.910 1.520 13.150 2.500 ;
        RECT  12.730 2.260 12.970 3.560 ;
        RECT  12.420 3.160 12.970 3.560 ;
        RECT  12.420 1.450 12.660 2.020 ;
        RECT  14.570 2.300 14.980 2.700 ;
        RECT  12.200 1.780 12.440 2.910 ;
        RECT  14.570 2.440 16.710 2.680 ;
        RECT  14.570 2.440 15.170 2.700 ;
        RECT  11.940 2.670 12.440 2.910 ;
        RECT  14.570 2.300 14.890 4.100 ;
        RECT  11.710 3.860 14.890 4.100 ;
        RECT  11.940 2.670 12.180 4.190 ;
        RECT  11.710 3.780 12.180 4.190 ;
        RECT  14.090 1.610 15.430 1.850 ;
        RECT  15.190 1.610 15.430 2.180 ;
        RECT  15.190 1.940 17.200 2.180 ;
        RECT  13.390 2.030 13.630 2.620 ;
        RECT  18.410 2.040 20.370 2.460 ;
        RECT  14.090 1.610 14.330 2.620 ;
        RECT  13.390 2.380 14.330 2.620 ;
        RECT  16.960 1.940 17.200 3.390 ;
        RECT  15.600 3.150 17.200 3.390 ;
        RECT  14.030 2.380 14.270 3.420 ;
        RECT  18.410 2.040 18.660 3.940 ;
        RECT  17.930 3.700 18.660 3.940 ;
        RECT  15.600 3.150 15.840 4.350 ;
        RECT  17.930 3.700 18.170 4.350 ;
        RECT  15.600 4.110 18.170 4.350 ;
    END
END mffnrb4

MACRO mffnrb2
    CLASS CORE ;
    FOREIGN mffnrb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.230  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.040 2.580 5.540 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.080 3.140 2.740 3.580 ;
        RECT  2.080 2.580 2.320 3.580 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.310 0.500 3.580 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.289  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.210 1.770 14.490 3.580 ;
        RECT  14.060 2.580 14.490 3.020 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.289  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.640 2.580 16.180 3.020 ;
        RECT  15.640 1.770 15.920 3.020 ;
        RECT  15.640 1.770 15.880 3.580 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  16.250 4.710 16.650 5.600 ;
        RECT  14.930 4.070 15.170 5.600 ;
        RECT  12.780 4.670 13.860 5.600 ;
        RECT  9.000 4.710 9.400 5.600 ;
        RECT  4.840 4.410 5.080 5.600 ;
        RECT  1.670 4.710 2.070 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  16.250 0.000 16.650 0.890 ;
        RECT  14.890 0.000 15.290 0.890 ;
        RECT  13.580 0.000 13.820 1.320 ;
        RECT  12.070 0.000 12.470 0.890 ;
        RECT  9.130 0.000 9.520 0.890 ;
        RECT  4.830 0.000 7.250 0.890 ;
        RECT  4.830 0.000 5.770 1.300 ;
        RECT  1.670 0.000 2.070 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.840 2.610 1.360 3.010 ;
        RECT  0.840 1.770 1.080 3.760 ;
        RECT  2.570 1.930 2.810 2.900 ;
        RECT  2.570 2.660 3.220 2.900 ;
        RECT  2.980 2.660 3.220 4.060 ;
        RECT  2.590 3.820 3.220 4.060 ;
        RECT  2.590 3.820 2.830 4.600 ;
        RECT  0.850 0.980 1.170 1.370 ;
        RECT  2.290 1.060 3.900 1.300 ;
        RECT  0.850 1.130 2.530 1.370 ;
        RECT  1.600 1.130 1.840 3.510 ;
        RECT  1.330 3.270 1.840 3.510 ;
        RECT  1.330 3.270 1.570 4.480 ;
        RECT  0.850 4.240 1.570 4.480 ;
        RECT  4.070 2.020 4.310 4.620 ;
        RECT  6.260 2.770 6.940 3.010 ;
        RECT  6.260 2.080 6.500 3.770 ;
        RECT  6.010 1.260 7.210 1.500 ;
        RECT  6.010 1.260 6.250 1.780 ;
        RECT  3.460 1.540 6.250 1.780 ;
        RECT  3.230 1.810 3.700 2.210 ;
        RECT  6.960 1.260 7.210 2.240 ;
        RECT  7.190 2.000 7.430 3.730 ;
        RECT  6.880 3.490 7.430 3.730 ;
        RECT  3.460 1.540 3.700 4.620 ;
        RECT  3.250 4.300 3.700 4.620 ;
        RECT  8.440 1.610 8.680 3.810 ;
        RECT  7.700 1.130 9.400 1.370 ;
        RECT  9.160 1.130 9.400 2.520 ;
        RECT  9.160 2.280 9.720 2.520 ;
        RECT  7.700 1.130 7.940 3.810 ;
        RECT  9.730 1.750 10.290 1.990 ;
        RECT  10.050 1.750 10.290 2.990 ;
        RECT  10.050 2.750 10.640 2.990 ;
        RECT  8.920 2.880 9.160 3.730 ;
        RECT  8.920 3.490 10.640 3.730 ;
        RECT  10.400 2.750 10.640 4.090 ;
        RECT  10.400 3.850 10.970 4.090 ;
        RECT  4.790 2.100 6.020 2.340 ;
        RECT  4.790 3.450 6.020 3.690 ;
        RECT  5.780 2.100 6.020 4.470 ;
        RECT  5.780 4.230 10.160 4.470 ;
        RECT  9.920 4.380 11.130 4.620 ;
        RECT  11.290 1.360 11.530 2.030 ;
        RECT  12.250 1.480 12.490 2.030 ;
        RECT  11.290 1.790 12.490 2.030 ;
        RECT  11.830 1.790 12.070 3.910 ;
        RECT  11.830 3.670 12.380 3.910 ;
        RECT  12.730 1.770 13.110 2.090 ;
        RECT  12.730 1.770 12.970 2.510 ;
        RECT  12.340 2.270 12.970 2.510 ;
        RECT  12.340 2.270 12.580 3.400 ;
        RECT  12.340 3.160 13.180 3.400 ;
        RECT  10.550 1.670 10.790 2.510 ;
        RECT  10.550 2.270 11.530 2.510 ;
        RECT  13.230 2.370 13.470 2.920 ;
        RECT  11.290 4.020 11.610 4.200 ;
        RECT  11.290 2.270 11.530 4.200 ;
        RECT  13.460 2.680 13.700 4.390 ;
        RECT  11.370 4.150 13.700 4.390 ;
    END
END mffnrb2

MACRO mffnrb1
    CLASS CORE ;
    FOREIGN mffnrb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.230  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.040 2.580 5.540 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.080 3.140 2.740 3.580 ;
        RECT  2.080 2.580 2.320 3.580 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.310 0.500 3.580 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.070 3.140 15.060 3.580 ;
        RECT  14.070 1.630 14.390 3.580 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.630 1.630 15.870 3.560 ;
        RECT  15.180 2.020 15.870 2.460 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  14.890 4.240 15.130 5.600 ;
        RECT  12.780 4.670 13.730 5.600 ;
        RECT  8.970 4.710 9.370 5.600 ;
        RECT  4.840 4.410 5.080 5.600 ;
        RECT  1.670 4.710 2.070 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  14.890 0.000 15.130 1.450 ;
        RECT  13.450 0.000 13.690 1.070 ;
        RECT  11.840 0.000 12.240 0.890 ;
        RECT  9.130 0.000 9.520 0.890 ;
        RECT  4.830 0.000 7.250 0.890 ;
        RECT  4.830 0.000 5.770 1.300 ;
        RECT  1.670 0.000 2.070 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.840 2.610 1.360 3.010 ;
        RECT  0.840 1.770 1.080 3.760 ;
        RECT  2.570 1.930 2.810 2.900 ;
        RECT  2.570 2.660 3.220 2.900 ;
        RECT  2.980 2.660 3.220 4.060 ;
        RECT  2.590 3.820 3.220 4.060 ;
        RECT  2.590 3.820 2.830 4.600 ;
        RECT  2.290 1.060 3.900 1.300 ;
        RECT  0.850 1.130 2.530 1.370 ;
        RECT  1.600 1.130 1.840 3.510 ;
        RECT  1.330 3.270 1.840 3.510 ;
        RECT  1.330 3.270 1.570 4.480 ;
        RECT  0.850 4.240 1.570 4.480 ;
        RECT  4.070 2.020 4.310 4.620 ;
        RECT  6.260 2.770 6.940 3.010 ;
        RECT  6.260 2.080 6.500 3.770 ;
        RECT  6.010 1.260 7.210 1.500 ;
        RECT  6.010 1.260 6.250 1.780 ;
        RECT  3.460 1.540 6.250 1.780 ;
        RECT  3.230 1.810 3.700 2.210 ;
        RECT  6.960 1.260 7.210 2.240 ;
        RECT  7.190 2.000 7.430 3.810 ;
        RECT  6.880 3.490 7.430 3.810 ;
        RECT  3.460 1.540 3.700 4.620 ;
        RECT  3.250 4.300 3.700 4.620 ;
        RECT  8.440 1.610 8.680 3.810 ;
        RECT  7.700 1.130 9.400 1.370 ;
        RECT  9.160 1.130 9.400 2.520 ;
        RECT  9.160 2.280 9.720 2.520 ;
        RECT  7.700 1.130 7.940 3.810 ;
        RECT  9.770 1.750 10.340 1.990 ;
        RECT  8.920 2.880 9.160 3.730 ;
        RECT  8.920 3.490 10.340 3.730 ;
        RECT  10.100 1.750 10.340 4.090 ;
        RECT  10.090 3.490 10.340 4.090 ;
        RECT  10.090 3.850 10.970 4.090 ;
        RECT  4.790 2.100 6.020 2.340 ;
        RECT  4.790 3.450 6.020 3.690 ;
        RECT  5.780 2.100 6.020 4.470 ;
        RECT  5.780 4.230 9.850 4.470 ;
        RECT  9.610 4.380 11.250 4.620 ;
        RECT  11.330 1.360 11.570 2.110 ;
        RECT  11.330 1.870 12.580 2.110 ;
        RECT  12.060 1.870 12.580 2.190 ;
        RECT  12.060 1.870 12.300 3.910 ;
        RECT  12.550 2.630 13.120 2.870 ;
        RECT  12.880 1.420 13.120 3.480 ;
        RECT  12.870 2.630 13.120 3.480 ;
        RECT  10.590 1.670 10.830 2.670 ;
        RECT  10.590 2.430 11.530 2.670 ;
        RECT  11.290 2.430 11.530 3.720 ;
        RECT  11.530 3.480 11.770 4.390 ;
        RECT  13.370 2.540 13.610 4.390 ;
        RECT  11.530 4.150 13.610 4.390 ;
    END
END mffnrb1

MACRO lanlq4
    CLASS CORE ;
    FOREIGN lanlq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.460 2.730 2.250 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.150 0.800 2.650 ;
        RECT  0.120 2.150 0.500 3.160 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.166  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.450 2.580 8.900 3.020 ;
        RECT  8.450 1.660 8.690 4.370 ;
        RECT  6.600 1.660 8.690 1.900 ;
        RECT  8.080 1.280 8.320 1.900 ;
        RECT  7.110 1.660 7.350 4.320 ;
        RECT  6.600 1.280 6.840 1.900 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  8.970 4.620 9.370 5.600 ;
        RECT  7.710 3.240 7.950 5.600 ;
        RECT  6.460 4.620 6.860 5.600 ;
        RECT  5.200 4.400 5.450 5.600 ;
        RECT  2.190 4.620 2.590 5.600 ;
        RECT  0.830 4.040 1.070 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.740 0.000 9.140 1.190 ;
        RECT  7.260 0.000 7.660 1.100 ;
        RECT  5.550 0.000 5.950 0.980 ;
        RECT  2.330 0.000 2.730 0.980 ;
        RECT  0.970 0.000 1.210 1.430 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.030 0.470 1.910 ;
        RECT  0.230 1.670 1.480 1.910 ;
        RECT  1.090 1.670 1.480 2.340 ;
        RECT  1.090 1.670 1.330 3.650 ;
        RECT  0.150 3.410 1.330 3.650 ;
        RECT  3.000 1.320 3.240 1.980 ;
        RECT  2.970 1.810 3.210 2.680 ;
        RECT  2.860 2.460 3.100 3.450 ;
        RECT  1.630 1.030 2.020 1.430 ;
        RECT  1.780 1.030 2.020 2.920 ;
        RECT  1.570 2.670 1.810 3.930 ;
        RECT  3.450 2.250 3.690 3.930 ;
        RECT  1.570 3.690 3.690 3.930 ;
        RECT  4.510 1.590 4.750 2.240 ;
        RECT  4.430 2.050 4.670 4.250 ;
        RECT  4.430 3.810 4.860 4.250 ;
        RECT  3.690 0.980 5.280 1.220 ;
        RECT  5.040 1.220 5.570 1.460 ;
        RECT  3.690 0.980 4.190 1.790 ;
        RECT  5.330 1.220 5.570 2.270 ;
        RECT  5.330 2.030 5.830 2.270 ;
        RECT  5.590 2.030 5.830 2.740 ;
        RECT  3.930 0.980 4.190 4.540 ;
        RECT  3.570 4.300 4.190 4.540 ;
        RECT  5.810 1.320 6.360 1.720 ;
        RECT  4.910 2.590 5.150 3.440 ;
        RECT  6.120 1.320 6.360 3.440 ;
        RECT  4.910 3.200 6.360 3.440 ;
    END
END lanlq4

MACRO lanlq2
    CLASS CORE ;
    FOREIGN lanlq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.401  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 2.580 2.740 3.020 ;
        RECT  2.220 2.580 2.550 3.460 ;
        RECT  2.220 1.940 2.460 3.460 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.500 3.490 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.200 3.140 7.780 3.580 ;
        RECT  7.200 1.770 7.440 3.580 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.820 4.070 8.060 5.600 ;
        RECT  6.500 4.070 6.740 5.600 ;
        RECT  4.900 4.710 5.300 5.600 ;
        RECT  2.150 4.240 2.390 5.600 ;
        RECT  0.610 4.390 0.850 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.870 0.000 8.110 1.600 ;
        RECT  6.460 0.000 6.700 1.590 ;
        RECT  5.010 0.000 5.250 1.440 ;
        RECT  2.040 0.000 2.280 1.250 ;
        RECT  0.480 0.000 0.880 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.420 1.310 0.980 1.550 ;
        RECT  0.740 1.310 0.980 3.970 ;
        RECT  0.420 3.730 0.980 3.970 ;
        RECT  1.260 2.450 1.830 2.690 ;
        RECT  1.260 1.410 1.500 3.990 ;
        RECT  1.260 3.670 1.700 3.990 ;
        RECT  2.660 1.490 3.250 1.730 ;
        RECT  3.010 1.490 3.250 4.020 ;
        RECT  2.710 3.700 3.250 4.020 ;
        RECT  4.260 1.410 4.510 3.990 ;
        RECT  3.520 1.410 3.770 4.470 ;
        RECT  5.260 2.770 5.500 4.470 ;
        RECT  3.520 4.230 5.500 4.470 ;
        RECT  4.750 2.020 6.000 2.260 ;
        RECT  5.760 1.410 6.000 3.990 ;
    END
END lanlq2

MACRO lanlq1
    CLASS CORE ;
    FOREIGN lanlq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.401  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 2.580 2.740 3.020 ;
        RECT  2.220 2.580 2.550 3.460 ;
        RECT  2.220 1.940 2.460 3.460 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.500 3.490 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.120 3.130 7.720 3.450 ;
        RECT  7.340 1.720 7.720 3.450 ;
        RECT  7.120 1.720 7.720 2.090 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  6.460 4.130 6.700 5.600 ;
        RECT  4.900 4.710 5.300 5.600 ;
        RECT  2.150 4.240 2.390 5.600 ;
        RECT  0.610 4.390 0.850 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.460 0.000 6.700 1.540 ;
        RECT  5.010 0.000 5.250 1.440 ;
        RECT  2.040 0.000 2.280 1.250 ;
        RECT  0.480 0.000 0.880 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.420 1.310 0.980 1.550 ;
        RECT  0.740 1.310 0.980 3.970 ;
        RECT  0.420 3.730 0.980 3.970 ;
        RECT  1.260 2.450 1.830 2.690 ;
        RECT  1.260 1.410 1.500 3.990 ;
        RECT  1.260 3.670 1.700 3.990 ;
        RECT  2.660 1.490 3.250 1.730 ;
        RECT  3.010 1.490 3.250 4.020 ;
        RECT  2.710 3.700 3.250 4.020 ;
        RECT  4.260 1.410 4.510 3.990 ;
        RECT  3.520 1.410 3.770 4.470 ;
        RECT  5.260 2.770 5.500 4.470 ;
        RECT  3.520 4.230 5.500 4.470 ;
        RECT  4.750 2.020 6.000 2.260 ;
        RECT  5.760 1.410 6.000 3.990 ;
    END
END lanlq1

MACRO lanln4
    CLASS CORE ;
    FOREIGN lanln4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.530 1.840 3.770 2.390 ;
        RECT  2.300 1.840 3.770 2.080 ;
        RECT  2.300 1.840 2.740 2.460 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.322  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 3.140 9.460 3.580 ;
        RECT  9.200 2.460 9.440 3.580 ;
        END
    END EN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.135  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.730 3.790 2.590 4.030 ;
        RECT  0.150 1.380 2.080 1.620 ;
        RECT  0.620 2.020 1.060 2.460 ;
        RECT  0.730 3.790 1.050 4.110 ;
        RECT  0.810 2.020 1.050 4.110 ;
        RECT  0.230 2.020 1.060 2.260 ;
        RECT  0.230 1.380 0.550 2.260 ;
        RECT  0.150 1.380 0.550 1.780 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  9.020 4.700 9.420 5.600 ;
        RECT  6.880 4.340 7.120 5.600 ;
        RECT  3.330 4.620 4.270 5.600 ;
        RECT  1.530 4.450 1.770 5.600 ;
        RECT  0.230 3.040 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  9.610 0.000 9.850 1.330 ;
        RECT  6.690 0.000 7.090 0.890 ;
        RECT  3.710 0.000 4.110 0.890 ;
        RECT  2.450 0.000 2.850 0.890 ;
        RECT  0.920 0.000 1.320 1.140 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.120 1.360 4.250 1.600 ;
        RECT  4.010 1.360 4.250 2.100 ;
        RECT  4.010 1.860 4.580 2.100 ;
        RECT  4.340 1.860 4.580 2.890 ;
        RECT  3.280 2.650 4.580 2.890 ;
        RECT  4.490 1.360 5.070 1.600 ;
        RECT  4.830 1.360 5.070 3.580 ;
        RECT  4.690 3.180 5.090 3.580 ;
        RECT  5.830 1.620 6.410 1.860 ;
        RECT  5.830 1.620 6.070 3.310 ;
        RECT  5.830 3.070 6.240 3.310 ;
        RECT  6.140 3.090 6.380 3.620 ;
        RECT  7.450 1.720 7.690 2.350 ;
        RECT  6.390 2.100 7.690 2.350 ;
        RECT  6.390 2.100 6.630 2.850 ;
        RECT  6.630 2.610 6.870 3.480 ;
        RECT  6.630 3.240 7.760 3.480 ;
        RECT  7.120 2.600 8.240 2.840 ;
        RECT  1.550 2.080 1.790 3.430 ;
        RECT  1.550 3.190 4.220 3.430 ;
        RECT  5.350 1.770 5.590 4.280 ;
        RECT  5.350 3.860 8.240 3.980 ;
        RECT  3.980 3.190 4.220 4.200 ;
        RECT  7.340 3.740 8.240 3.980 ;
        RECT  8.000 2.600 8.240 3.980 ;
        RECT  3.980 3.950 7.580 4.100 ;
        RECT  3.980 3.950 5.690 4.200 ;
        RECT  5.290 3.870 5.690 4.280 ;
        RECT  5.630 1.050 6.420 1.290 ;
        RECT  6.190 1.130 8.170 1.370 ;
        RECT  7.930 1.130 8.170 1.990 ;
        RECT  7.930 1.750 8.780 1.990 ;
        RECT  8.520 1.750 8.780 4.540 ;
        RECT  8.070 4.300 8.780 4.540 ;
        RECT  8.410 1.050 9.370 1.290 ;
        RECT  9.130 1.050 9.370 2.040 ;
        RECT  9.130 1.720 9.960 2.040 ;
        RECT  9.540 1.720 9.960 2.120 ;
        RECT  9.720 1.720 9.960 4.310 ;
        RECT  9.530 3.850 9.960 4.310 ;
    END
END lanln4

MACRO lanln2
    CLASS CORE ;
    FOREIGN lanln2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.020 2.740 2.460 ;
        RECT  2.300 2.020 2.700 3.540 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.960 ;
        END
    END EN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.400 3.140 8.900 3.580 ;
        RECT  8.400 1.770 8.640 3.580 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  9.020 4.070 9.260 5.600 ;
        RECT  7.700 4.070 7.940 5.600 ;
        RECT  6.330 4.430 6.570 5.600 ;
        RECT  3.640 3.930 3.880 5.600 ;
        RECT  2.200 3.960 2.440 5.600 ;
        RECT  0.630 3.830 0.870 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.970 0.000 9.370 0.990 ;
        RECT  7.550 0.000 7.940 1.080 ;
        RECT  6.430 0.000 6.820 1.030 ;
        RECT  3.490 0.000 3.730 1.200 ;
        RECT  2.100 0.000 2.500 1.090 ;
        RECT  0.580 0.000 0.980 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.630 1.230 0.980 1.550 ;
        RECT  0.740 2.050 1.250 2.450 ;
        RECT  0.740 1.230 0.980 3.490 ;
        RECT  0.630 3.170 0.980 3.490 ;
        RECT  1.330 1.490 1.740 1.810 ;
        RECT  1.490 2.460 2.050 2.860 ;
        RECT  1.490 1.490 1.740 4.260 ;
        RECT  1.380 3.940 1.740 4.260 ;
        RECT  2.710 1.540 4.020 1.780 ;
        RECT  3.690 1.540 4.020 1.980 ;
        RECT  3.690 1.540 3.930 3.340 ;
        RECT  2.940 3.100 3.930 3.340 ;
        RECT  2.940 3.100 3.180 4.260 ;
        RECT  4.260 1.130 4.500 3.710 ;
        RECT  5.620 1.430 6.060 1.750 ;
        RECT  5.620 1.430 5.860 3.710 ;
        RECT  5.620 3.390 6.060 3.710 ;
        RECT  6.300 2.600 7.180 2.840 ;
        RECT  5.000 1.430 5.240 4.190 ;
        RECT  6.300 2.600 6.540 4.190 ;
        RECT  5.000 3.950 6.540 4.190 ;
        RECT  7.110 1.430 7.350 2.280 ;
        RECT  6.100 2.040 7.670 2.280 ;
        RECT  7.430 2.040 7.670 3.630 ;
        RECT  7.030 3.390 7.670 3.630 ;
    END
END lanln2

MACRO lanln1
    CLASS CORE ;
    FOREIGN lanln1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.020 2.740 2.460 ;
        RECT  2.300 2.020 2.700 3.540 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.960 ;
        END
    END EN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 1.430 8.840 3.450 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.750 4.130 7.990 5.600 ;
        RECT  6.330 4.430 6.570 5.600 ;
        RECT  3.640 3.930 3.880 5.600 ;
        RECT  2.200 3.960 2.440 5.600 ;
        RECT  0.630 3.830 0.870 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.630 0.000 8.040 1.070 ;
        RECT  6.480 0.000 6.720 1.770 ;
        RECT  3.490 0.000 3.730 1.200 ;
        RECT  2.100 0.000 2.500 1.090 ;
        RECT  0.580 0.000 0.980 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.630 1.230 0.980 1.550 ;
        RECT  0.740 2.040 1.250 2.440 ;
        RECT  0.740 1.230 0.980 3.490 ;
        RECT  0.630 3.170 0.980 3.490 ;
        RECT  1.330 1.490 1.740 1.810 ;
        RECT  1.490 2.460 2.050 2.860 ;
        RECT  1.490 1.490 1.740 4.260 ;
        RECT  1.380 3.940 1.740 4.260 ;
        RECT  2.710 1.540 4.020 1.780 ;
        RECT  3.690 1.540 4.020 1.980 ;
        RECT  3.690 1.540 3.930 3.340 ;
        RECT  2.940 3.100 3.930 3.340 ;
        RECT  2.940 3.100 3.180 4.260 ;
        RECT  4.260 1.130 4.500 3.710 ;
        RECT  5.700 1.430 6.060 1.750 ;
        RECT  5.700 1.430 5.940 3.710 ;
        RECT  5.700 3.390 6.060 3.710 ;
        RECT  6.300 2.850 7.180 3.090 ;
        RECT  5.000 1.430 5.240 4.190 ;
        RECT  6.300 2.850 6.540 4.190 ;
        RECT  5.000 3.950 6.540 4.190 ;
        RECT  7.220 1.430 7.460 2.280 ;
        RECT  6.180 2.040 7.670 2.280 ;
        RECT  7.430 2.040 7.670 3.630 ;
        RECT  7.030 3.390 7.670 3.630 ;
    END
END lanln1

MACRO lanlb4
    CLASS CORE ;
    FOREIGN lanlb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 1.570 4.590 2.170 ;
        RECT  3.980 1.460 4.420 2.170 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.820 2.300 12.200 3.020 ;
        RECT  11.460 2.300 12.200 2.540 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.689  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.150 3.370 3.230 3.610 ;
        RECT  1.560 1.540 2.100 1.800 ;
        RECT  0.160 1.640 1.770 1.880 ;
        RECT  0.120 2.540 0.560 3.370 ;
        RECT  0.320 1.540 0.560 3.610 ;
        RECT  0.150 2.540 0.550 3.690 ;
        RECT  0.160 1.540 0.560 1.940 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.987  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.400 1.600 9.970 1.840 ;
        RECT  7.520 1.610 9.480 1.850 ;
        RECT  8.880 2.580 9.460 3.240 ;
        RECT  7.520 2.920 9.460 3.160 ;
        RECT  8.870 2.580 9.460 3.160 ;
        RECT  7.520 1.610 7.920 3.230 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.320 5.600 ;
        RECT  11.000 4.490 11.400 5.600 ;
        RECT  9.560 4.400 9.960 5.600 ;
        RECT  8.260 4.400 8.660 5.600 ;
        RECT  6.960 4.400 7.360 5.600 ;
        RECT  4.160 4.710 4.560 5.600 ;
        RECT  2.240 3.950 2.640 5.600 ;
        RECT  0.780 4.020 1.180 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.320 0.740 ;
        RECT  11.030 0.000 11.430 1.000 ;
        RECT  8.790 0.000 9.190 0.890 ;
        RECT  7.250 0.000 7.650 0.890 ;
        RECT  2.470 0.000 3.410 0.890 ;
        RECT  0.930 0.000 1.330 1.330 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  4.620 1.080 5.200 1.320 ;
        RECT  4.960 1.080 5.200 2.410 ;
        RECT  4.910 2.140 5.150 3.460 ;
        RECT  3.240 2.410 4.330 2.650 ;
        RECT  4.090 2.410 4.330 3.960 ;
        RECT  5.440 1.000 5.680 3.960 ;
        RECT  4.090 3.720 5.900 3.960 ;
        RECT  5.510 3.640 5.900 4.040 ;
        RECT  6.410 1.520 6.650 3.450 ;
        RECT  6.170 3.050 6.650 3.450 ;
        RECT  2.760 1.520 3.470 1.760 ;
        RECT  2.760 1.520 3.000 3.130 ;
        RECT  2.760 2.890 3.850 3.130 ;
        RECT  6.890 2.190 7.130 4.160 ;
        RECT  6.390 3.920 7.130 4.160 ;
        RECT  3.610 2.890 3.850 4.440 ;
        RECT  3.610 4.200 5.200 4.440 ;
        RECT  6.390 3.920 6.630 4.520 ;
        RECT  5.010 4.280 6.630 4.520 ;
        RECT  5.920 1.040 7.030 1.280 ;
        RECT  9.260 1.120 10.580 1.360 ;
        RECT  6.840 1.130 9.330 1.370 ;
        RECT  5.920 1.040 6.160 2.610 ;
        RECT  10.340 1.120 10.580 3.630 ;
        RECT  10.830 1.600 12.120 1.840 ;
        RECT  10.830 1.600 11.070 3.550 ;
        RECT  10.830 3.310 12.170 3.550 ;
    END
END lanlb4

MACRO lanlb2
    CLASS CORE ;
    FOREIGN lanlb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.337  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.460 2.900 3.410 ;
        RECT  2.300 1.460 2.900 1.900 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.254  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.340 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 1.370 7.670 1.700 ;
        RECT  7.290 1.370 7.530 3.740 ;
        RECT  6.780 1.370 7.530 1.900 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 3.140 8.990 3.740 ;
        RECT  8.750 1.380 8.990 3.740 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  9.300 4.290 9.540 5.600 ;
        RECT  7.880 4.290 8.120 5.600 ;
        RECT  6.580 4.290 6.820 5.600 ;
        RECT  5.210 4.690 5.610 5.600 ;
        RECT  2.300 4.050 2.540 5.600 ;
        RECT  0.500 4.490 0.740 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  9.470 0.000 9.710 1.260 ;
        RECT  8.050 0.000 8.290 1.240 ;
        RECT  6.570 0.000 6.970 0.970 ;
        RECT  5.130 0.000 5.530 0.890 ;
        RECT  2.400 0.000 2.640 1.220 ;
        RECT  0.630 0.000 1.030 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.840 1.230 1.320 1.550 ;
        RECT  1.080 1.230 1.320 4.070 ;
        RECT  0.570 3.830 1.320 4.070 ;
        RECT  1.560 2.410 2.290 2.650 ;
        RECT  1.560 1.000 1.900 3.750 ;
        RECT  3.140 1.360 3.380 3.980 ;
        RECT  2.960 3.660 3.380 3.980 ;
        RECT  4.620 1.350 4.860 2.020 ;
        RECT  4.520 1.780 4.760 3.940 ;
        RECT  5.000 2.940 5.870 3.180 ;
        RECT  3.880 1.360 4.120 4.420 ;
        RECT  3.780 3.540 4.120 4.420 ;
        RECT  5.000 2.940 5.240 4.420 ;
        RECT  3.780 4.180 5.240 4.420 ;
        RECT  5.980 1.360 6.220 2.700 ;
        RECT  5.000 2.260 6.220 2.500 ;
        RECT  5.980 2.460 7.050 2.700 ;
        RECT  6.110 2.460 6.350 3.860 ;
        RECT  5.800 3.620 6.350 3.860 ;
    END
END lanlb2

MACRO lanlb1
    CLASS CORE ;
    FOREIGN lanlb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.337  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.890 3.090 2.290 ;
        RECT  2.650 1.890 2.900 3.410 ;
        RECT  2.300 1.460 2.740 2.130 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.254  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.340 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.973  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.530 1.420 7.220 1.900 ;
        RECT  6.790 1.420 7.030 3.320 ;
        RECT  6.580 3.080 6.820 3.740 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.995  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.880 2.580 8.170 3.740 ;
        RECT  7.930 1.420 8.170 3.740 ;
        RECT  7.340 2.580 8.170 3.020 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.170 4.360 7.410 5.600 ;
        RECT  5.210 4.660 5.610 5.600 ;
        RECT  2.300 4.050 2.540 5.600 ;
        RECT  0.500 4.490 0.740 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.190 0.000 7.590 1.180 ;
        RECT  5.060 0.000 5.460 0.890 ;
        RECT  2.150 0.000 2.570 0.890 ;
        RECT  0.630 0.000 1.030 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.840 1.230 1.320 1.550 ;
        RECT  1.080 1.230 1.320 4.070 ;
        RECT  0.570 3.830 1.320 4.070 ;
        RECT  1.560 2.490 2.290 2.730 ;
        RECT  1.560 1.360 1.900 3.940 ;
        RECT  2.990 1.410 3.570 1.650 ;
        RECT  3.330 1.410 3.570 3.080 ;
        RECT  3.270 2.840 3.510 3.900 ;
        RECT  2.960 3.660 3.510 3.900 ;
        RECT  4.550 1.350 4.790 2.020 ;
        RECT  4.520 1.780 4.760 3.940 ;
        RECT  5.000 3.030 5.860 3.270 ;
        RECT  3.810 1.360 4.050 4.420 ;
        RECT  3.780 3.540 4.050 4.420 ;
        RECT  5.000 3.030 5.240 4.420 ;
        RECT  3.780 4.180 5.240 4.420 ;
        RECT  5.910 1.340 6.150 2.590 ;
        RECT  5.000 2.350 6.550 2.590 ;
        RECT  6.100 2.350 6.550 2.700 ;
        RECT  6.100 2.350 6.340 3.940 ;
        RECT  5.800 3.620 6.340 3.940 ;
    END
END lanlb1

MACRO lanht4
    CLASS CORE ;
    FOREIGN lanht4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.280 2.580 2.740 3.040 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.322  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.990 0.540 2.390 ;
        RECT  0.120 2.580 0.500 3.020 ;
        RECT  0.140 1.990 0.500 3.020 ;
        END
    END E
    PIN OE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.886  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.580 2.580 10.260 3.020 ;
        RECT  10.020 2.040 10.260 3.020 ;
        END
    END OE
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.589  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.820 2.020 12.200 2.460 ;
        RECT  11.270 2.770 12.060 3.010 ;
        RECT  11.820 1.690 12.060 3.010 ;
        RECT  11.030 1.690 12.060 1.930 ;
        RECT  11.190 3.940 11.590 4.340 ;
        RECT  9.890 3.830 11.510 4.070 ;
        RECT  11.270 2.770 11.510 4.340 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.320 5.600 ;
        RECT  11.770 3.250 12.170 3.650 ;
        RECT  11.850 3.250 12.090 5.600 ;
        RECT  10.630 4.620 11.030 5.600 ;
        RECT  9.300 4.400 9.700 5.600 ;
        RECT  7.290 4.330 7.690 5.600 ;
        RECT  4.710 4.330 5.110 5.600 ;
        RECT  2.190 4.700 2.590 5.600 ;
        RECT  0.890 4.180 1.290 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.320 0.740 ;
        RECT  11.770 0.000 12.170 0.980 ;
        RECT  10.290 0.000 10.690 0.980 ;
        RECT  7.110 0.000 7.510 1.640 ;
        RECT  4.880 0.000 5.280 0.890 ;
        RECT  2.210 0.000 2.610 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.230 0.550 1.750 ;
        RECT  0.150 1.510 1.140 1.750 ;
        RECT  0.900 1.510 1.140 3.500 ;
        RECT  0.230 3.260 1.140 3.500 ;
        RECT  0.230 3.260 0.470 4.580 ;
        RECT  2.460 1.620 3.200 1.860 ;
        RECT  2.460 1.620 2.700 2.340 ;
        RECT  2.460 2.100 3.220 2.340 ;
        RECT  2.980 2.100 3.220 4.360 ;
        RECT  2.780 3.960 3.220 4.360 ;
        RECT  2.990 0.980 3.390 1.380 ;
        RECT  1.510 1.140 3.390 1.380 ;
        RECT  1.510 1.060 1.910 1.460 ;
        RECT  1.570 1.060 1.810 3.830 ;
        RECT  4.110 1.620 4.690 1.860 ;
        RECT  4.110 1.620 4.350 2.580 ;
        RECT  3.940 2.340 4.180 3.970 ;
        RECT  3.940 3.730 4.550 3.970 ;
        RECT  3.630 0.980 4.570 1.220 ;
        RECT  4.340 1.130 5.260 1.370 ;
        RECT  3.630 0.980 3.870 2.100 ;
        RECT  5.020 1.130 5.260 2.370 ;
        RECT  5.020 2.130 5.550 2.370 ;
        RECT  5.310 2.130 5.550 2.850 ;
        RECT  3.460 1.860 3.700 3.470 ;
        RECT  5.650 1.500 6.050 1.900 ;
        RECT  4.590 2.520 4.830 3.330 ;
        RECT  5.810 1.500 6.050 3.330 ;
        RECT  4.590 3.090 6.050 3.330 ;
        RECT  5.530 3.090 5.770 3.920 ;
        RECT  5.840 1.010 6.560 1.250 ;
        RECT  6.320 1.240 6.770 1.640 ;
        RECT  7.930 1.240 8.170 2.060 ;
        RECT  7.670 1.820 8.170 2.060 ;
        RECT  7.670 1.820 7.910 2.470 ;
        RECT  6.320 2.230 7.910 2.470 ;
        RECT  6.320 1.010 6.560 4.110 ;
        RECT  6.060 3.870 6.560 4.110 ;
        RECT  6.060 3.870 6.300 4.620 ;
        RECT  9.150 0.980 9.650 1.380 ;
        RECT  9.410 0.980 9.650 2.320 ;
        RECT  8.890 2.080 9.650 2.320 ;
        RECT  8.890 2.080 9.130 3.020 ;
        RECT  8.640 2.780 9.130 3.020 ;
        RECT  8.640 2.780 8.880 3.660 ;
        RECT  8.410 1.590 8.990 1.830 ;
        RECT  8.410 1.590 8.650 2.540 ;
        RECT  8.150 2.300 8.650 2.540 ;
        RECT  8.150 2.300 8.390 3.030 ;
        RECT  6.800 2.790 8.390 3.030 ;
        RECT  10.790 2.520 11.030 3.500 ;
        RECT  9.200 3.260 11.030 3.500 ;
        RECT  6.800 3.440 8.350 3.680 ;
        RECT  6.800 2.790 7.040 4.060 ;
        RECT  9.200 3.260 9.440 4.160 ;
        RECT  8.110 3.920 9.440 4.160 ;
        RECT  8.110 3.440 8.350 4.620 ;
    END
END lanht4

MACRO lanht2
    CLASS CORE ;
    FOREIGN lanht2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.410 1.420 2.650 ;
        RECT  0.620 2.020 1.060 2.650 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.890 0.500 3.580 ;
        END
    END E
    PIN OE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.758  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.990 2.260 7.810 2.500 ;
        RECT  6.780 2.020 7.220 2.500 ;
        END
    END OE
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.950 3.700 9.960 3.940 ;
        RECT  9.580 1.620 9.960 3.940 ;
        RECT  9.130 1.620 9.960 1.860 ;
        RECT  9.130 1.010 9.370 1.860 ;
        RECT  8.330 1.010 9.370 1.250 ;
        RECT  5.950 2.740 6.190 4.310 ;
        RECT  5.510 1.720 6.120 1.960 ;
        RECT  5.510 2.740 6.190 2.980 ;
        RECT  5.510 1.720 5.750 2.980 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  9.610 4.220 9.850 5.600 ;
        RECT  7.100 4.620 7.500 5.600 ;
        RECT  4.690 4.620 5.090 5.600 ;
        RECT  0.230 3.840 1.390 4.080 ;
        RECT  1.150 3.510 1.390 4.080 ;
        RECT  0.230 3.840 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  9.610 0.000 9.850 1.260 ;
        RECT  7.000 0.000 7.240 1.460 ;
        RECT  3.820 0.000 4.760 1.180 ;
        RECT  1.320 0.000 1.560 1.280 ;
        RECT  0.420 0.000 0.820 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.140 1.720 2.380 3.540 ;
        RECT  0.580 1.230 0.820 1.780 ;
        RECT  0.580 1.540 1.900 1.780 ;
        RECT  1.660 1.540 1.900 4.560 ;
        RECT  0.890 4.320 2.440 4.560 ;
        RECT  3.660 1.880 4.220 2.120 ;
        RECT  3.660 1.880 3.900 3.460 ;
        RECT  3.660 3.220 4.220 3.460 ;
        RECT  2.550 0.980 3.480 1.220 ;
        RECT  2.550 0.980 2.920 1.410 ;
        RECT  2.680 0.980 2.920 4.620 ;
        RECT  2.680 4.380 4.260 4.620 ;
        RECT  3.160 1.800 3.400 4.090 ;
        RECT  3.160 3.850 5.470 4.090 ;
        RECT  5.030 0.980 5.590 1.220 ;
        RECT  4.140 2.410 5.270 2.650 ;
        RECT  5.030 0.980 5.270 3.460 ;
        RECT  5.030 3.220 5.710 3.460 ;
        RECT  7.660 1.660 8.370 1.900 ;
        RECT  8.130 2.690 8.980 2.930 ;
        RECT  8.130 1.660 8.370 3.460 ;
        RECT  7.630 3.220 8.370 3.460 ;
    END
END lanht2

MACRO lanht1
    CLASS CORE ;
    FOREIGN lanht1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.410 1.420 2.650 ;
        RECT  0.620 2.020 1.060 2.650 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.890 0.500 3.580 ;
        END
    END E
    PIN OE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.441  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.900 2.180 8.280 3.020 ;
        RECT  7.600 2.180 8.280 2.500 ;
        END
    END OE
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.071  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.950 2.580 6.660 3.020 ;
        RECT  5.950 1.110 6.190 4.310 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.150 4.220 7.390 5.600 ;
        RECT  4.690 4.620 5.090 5.600 ;
        RECT  0.230 3.840 1.390 4.080 ;
        RECT  1.150 3.510 1.390 4.080 ;
        RECT  0.230 3.840 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.150 0.000 7.390 1.260 ;
        RECT  4.620 0.000 4.860 1.440 ;
        RECT  3.900 0.000 4.140 1.180 ;
        RECT  1.320 0.000 1.560 1.280 ;
        RECT  0.420 0.000 0.820 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.140 1.720 2.380 3.540 ;
        RECT  0.580 1.230 0.820 1.780 ;
        RECT  0.580 1.540 1.900 1.780 ;
        RECT  1.660 1.540 1.900 4.560 ;
        RECT  0.890 4.320 2.440 4.560 ;
        RECT  3.900 1.800 4.140 3.540 ;
        RECT  2.550 0.980 3.480 1.220 ;
        RECT  2.550 0.980 2.920 1.410 ;
        RECT  2.680 0.980 2.920 4.620 ;
        RECT  2.680 4.380 4.260 4.620 ;
        RECT  3.160 1.800 3.400 4.090 ;
        RECT  3.160 3.850 5.470 4.090 ;
        RECT  4.380 2.410 5.630 2.650 ;
        RECT  5.390 1.800 5.630 3.540 ;
        RECT  6.900 1.520 8.240 1.760 ;
        RECT  6.900 1.520 7.140 3.500 ;
        RECT  6.900 3.260 8.250 3.500 ;
    END
END lanht1

MACRO lanhq4
    CLASS CORE ;
    FOREIGN lanhq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.580 1.760 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.800 4.420 3.580 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.171  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.980 1.960 8.730 2.200 ;
        RECT  8.490 1.070 8.730 2.200 ;
        RECT  7.900 1.960 8.340 2.460 ;
        RECT  5.760 3.650 8.250 3.890 ;
        RECT  8.010 1.960 8.250 3.890 ;
        RECT  6.980 1.070 7.220 2.200 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.810 4.620 8.210 5.600 ;
        RECT  6.500 4.610 6.900 5.600 ;
        RECT  3.740 4.550 4.140 5.600 ;
        RECT  0.750 4.620 1.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.650 0.000 8.050 0.980 ;
        RECT  6.150 0.000 6.550 0.980 ;
        RECT  3.970 0.000 4.210 1.120 ;
        RECT  1.150 0.000 1.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.700 2.020 2.250 2.260 ;
        RECT  2.010 2.020 2.250 3.620 ;
        RECT  1.520 3.380 2.250 3.620 ;
        RECT  1.190 1.530 2.600 1.770 ;
        RECT  0.120 1.630 1.470 1.870 ;
        RECT  0.120 1.630 0.550 2.030 ;
        RECT  0.120 1.630 0.360 4.050 ;
        RECT  0.120 3.650 0.550 4.050 ;
        RECT  3.320 1.840 3.560 3.070 ;
        RECT  3.070 2.830 3.560 3.070 ;
        RECT  3.070 2.830 3.310 3.810 ;
        RECT  4.480 2.100 4.900 2.500 ;
        RECT  0.600 3.170 0.990 3.410 ;
        RECT  0.600 2.270 0.840 3.410 ;
        RECT  0.790 3.210 1.030 4.380 ;
        RECT  4.660 2.100 4.900 4.310 ;
        RECT  3.260 4.070 4.900 4.310 ;
        RECT  0.790 4.140 1.790 4.380 ;
        RECT  3.260 4.070 3.500 4.620 ;
        RECT  1.550 4.380 3.500 4.620 ;
        RECT  2.530 0.980 3.720 1.220 ;
        RECT  3.480 0.980 3.720 1.600 ;
        RECT  3.480 1.360 4.130 1.600 ;
        RECT  3.890 1.360 4.130 1.860 ;
        RECT  2.870 0.980 3.110 1.620 ;
        RECT  3.890 1.620 5.320 1.860 ;
        RECT  5.100 1.720 6.250 1.960 ;
        RECT  5.300 1.720 6.250 2.120 ;
        RECT  2.840 1.460 3.080 2.530 ;
        RECT  2.590 2.290 3.080 2.530 ;
        RECT  2.590 2.290 2.830 4.140 ;
        RECT  2.240 3.900 2.830 4.140 ;
        RECT  5.380 0.980 5.780 1.380 ;
        RECT  5.510 1.220 6.730 1.460 ;
        RECT  6.490 1.220 6.730 2.730 ;
        RECT  5.280 2.490 6.730 2.730 ;
        RECT  5.280 2.490 5.520 4.600 ;
        RECT  8.490 3.800 8.730 4.370 ;
        RECT  5.280 4.130 8.730 4.370 ;
        RECT  5.280 4.130 5.800 4.600 ;
    END
END lanhq4

MACRO lanhq2
    CLASS CORE ;
    FOREIGN lanhq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.306  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.500 1.960 2.740 3.480 ;
        RECT  2.260 1.960 2.740 2.460 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.540 3.380 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.248  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.080 3.140 7.780 3.580 ;
        RECT  7.540 1.850 7.780 3.580 ;
        RECT  7.140 1.850 7.780 2.090 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.870 4.070 8.110 5.600 ;
        RECT  6.570 4.070 6.810 5.600 ;
        RECT  5.510 4.180 5.750 5.600 ;
        RECT  2.250 3.870 2.490 5.600 ;
        RECT  0.640 4.280 0.880 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.930 0.000 8.170 1.620 ;
        RECT  6.530 0.000 6.770 1.620 ;
        RECT  5.050 0.000 5.290 1.370 ;
        RECT  2.090 0.000 2.330 1.710 ;
        RECT  0.530 0.000 0.770 1.430 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.530 1.850 1.110 2.090 ;
        RECT  0.870 1.850 1.110 3.860 ;
        RECT  0.460 3.620 1.110 3.860 ;
        RECT  1.270 1.390 1.840 1.630 ;
        RECT  1.600 1.390 1.840 4.010 ;
        RECT  1.430 3.690 1.840 4.010 ;
        RECT  2.750 1.400 3.230 1.720 ;
        RECT  2.990 1.400 3.230 4.010 ;
        RECT  4.230 1.430 4.570 1.750 ;
        RECT  4.330 1.430 4.570 4.010 ;
        RECT  4.330 3.690 4.790 4.010 ;
        RECT  3.490 1.430 3.970 1.750 ;
        RECT  5.030 2.600 5.900 2.840 ;
        RECT  3.730 1.430 3.970 4.490 ;
        RECT  5.030 2.600 5.270 4.490 ;
        RECT  3.730 4.250 5.270 4.490 ;
        RECT  5.830 1.430 6.070 2.280 ;
        RECT  4.810 2.040 6.380 2.280 ;
        RECT  6.140 2.040 6.380 3.660 ;
        RECT  5.750 3.420 6.380 3.660 ;
    END
END lanhq2

MACRO lanhq1
    CLASS CORE ;
    FOREIGN lanhq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.306  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.500 1.960 2.740 3.480 ;
        RECT  2.260 1.960 2.740 2.460 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.540 3.380 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.230  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.310 1.550 7.720 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  6.530 4.140 6.770 5.600 ;
        RECT  5.510 4.180 5.750 5.600 ;
        RECT  2.250 3.870 2.490 5.600 ;
        RECT  0.640 4.280 0.880 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.570 0.000 6.810 1.370 ;
        RECT  5.050 0.000 5.290 1.370 ;
        RECT  2.090 0.000 2.330 1.710 ;
        RECT  0.530 0.000 0.770 1.430 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.530 1.850 1.110 2.090 ;
        RECT  0.870 1.850 1.110 3.860 ;
        RECT  0.460 3.620 1.110 3.860 ;
        RECT  1.270 1.390 1.840 1.630 ;
        RECT  1.600 1.390 1.840 4.010 ;
        RECT  1.430 3.690 1.840 4.010 ;
        RECT  2.750 1.400 3.230 1.720 ;
        RECT  2.990 1.400 3.230 4.010 ;
        RECT  4.230 1.430 4.570 1.750 ;
        RECT  4.330 1.430 4.570 4.010 ;
        RECT  4.330 3.690 4.790 4.010 ;
        RECT  3.490 1.430 3.970 1.750 ;
        RECT  5.030 2.600 5.900 2.840 ;
        RECT  3.730 1.430 3.970 4.490 ;
        RECT  5.030 2.600 5.270 4.490 ;
        RECT  3.730 4.250 5.270 4.490 ;
        RECT  5.830 1.430 6.070 2.280 ;
        RECT  4.810 2.040 6.380 2.280 ;
        RECT  6.140 2.040 6.380 3.660 ;
        RECT  5.750 3.420 6.380 3.660 ;
    END
END lanhq1

MACRO lanhn4
    CLASS CORE ;
    FOREIGN lanhn4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.271  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.100 2.780 2.500 ;
        RECT  2.300 2.020 2.740 2.500 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.329  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.860 0.790 2.260 ;
        RECT  0.120 1.860 0.500 2.460 ;
        END
    END E
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.608  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 3.680 9.930 3.920 ;
        RECT  6.820 3.420 9.460 3.820 ;
        RECT  9.020 1.120 9.460 3.920 ;
        RECT  8.670 1.090 9.390 1.480 ;
        RECT  8.950 1.120 9.460 1.520 ;
        RECT  7.500 1.230 9.460 1.480 ;
        RECT  7.160 1.170 7.740 1.410 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  8.860 4.610 9.260 5.600 ;
        RECT  7.380 4.170 7.780 5.600 ;
        RECT  5.520 4.400 5.920 5.600 ;
        RECT  2.090 4.710 2.490 5.600 ;
        RECT  0.740 4.680 1.140 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  9.530 0.000 9.930 0.890 ;
        RECT  7.920 0.000 8.320 0.990 ;
        RECT  5.690 0.000 6.090 0.890 ;
        RECT  2.660 0.000 3.060 0.890 ;
        RECT  0.730 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.380 1.270 1.620 ;
        RECT  1.030 1.380 1.270 2.740 ;
        RECT  1.030 1.840 1.480 2.240 ;
        RECT  0.740 2.500 1.280 2.740 ;
        RECT  1.030 1.840 1.280 2.740 ;
        RECT  0.480 2.700 0.980 2.940 ;
        RECT  0.480 2.700 0.720 4.250 ;
        RECT  0.150 4.010 0.720 4.250 ;
        RECT  2.210 1.540 3.430 1.780 ;
        RECT  3.190 1.540 3.430 2.800 ;
        RECT  3.060 2.400 3.460 2.800 ;
        RECT  3.020 2.530 3.260 3.190 ;
        RECT  2.040 2.950 3.260 3.190 ;
        RECT  3.670 1.020 3.910 2.100 ;
        RECT  3.710 1.850 3.950 3.220 ;
        RECT  3.650 2.970 3.890 4.050 ;
        RECT  3.300 3.810 3.890 4.050 ;
        RECT  1.510 1.000 2.440 1.240 ;
        RECT  1.510 1.000 1.960 1.560 ;
        RECT  1.720 1.000 1.960 2.720 ;
        RECT  1.520 2.480 1.760 3.440 ;
        RECT  1.340 3.040 1.760 3.440 ;
        RECT  1.420 2.940 1.660 4.470 ;
        RECT  1.420 4.230 3.020 4.470 ;
        RECT  2.780 4.380 4.820 4.620 ;
        RECT  4.810 1.610 5.510 1.850 ;
        RECT  4.810 1.610 5.050 3.530 ;
        RECT  4.190 1.020 4.730 1.370 ;
        RECT  4.190 1.130 6.300 1.370 ;
        RECT  4.190 1.020 4.660 1.420 ;
        RECT  6.060 1.130 6.300 2.600 ;
        RECT  6.060 2.200 8.300 2.600 ;
        RECT  4.190 1.020 4.430 3.720 ;
        RECT  4.140 3.480 4.380 4.120 ;
        RECT  6.540 0.980 6.780 1.960 ;
        RECT  6.540 1.720 8.780 1.960 ;
        RECT  5.350 2.230 5.590 3.130 ;
        RECT  8.540 1.720 8.780 3.130 ;
        RECT  5.350 2.890 8.780 3.130 ;
        RECT  6.200 2.890 6.440 3.740 ;
    END
END lanhn4

MACRO lanhn2
    CLASS CORE ;
    FOREIGN lanhn2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.700 2.740 4.200 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.480 ;
        END
    END E
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.310 1.460 8.900 2.490 ;
        RECT  8.310 1.110 8.550 3.450 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  9.050 4.130 9.290 5.600 ;
        RECT  7.460 4.470 7.860 5.600 ;
        RECT  6.460 4.710 6.860 5.600 ;
        RECT  3.300 3.840 3.540 5.600 ;
        RECT  1.780 3.700 2.020 5.600 ;
        RECT  0.420 4.710 0.820 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.970 0.000 9.370 0.980 ;
        RECT  7.460 0.000 7.860 0.980 ;
        RECT  6.300 0.000 6.540 1.550 ;
        RECT  3.310 0.000 3.550 1.200 ;
        RECT  2.220 0.000 2.460 1.200 ;
        RECT  0.720 0.000 0.960 1.210 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 2.600 1.760 2.840 ;
        RECT  0.740 1.550 0.980 2.960 ;
        RECT  0.440 2.720 0.980 2.960 ;
        RECT  0.440 2.720 0.680 4.370 ;
        RECT  0.440 4.050 0.820 4.370 ;
        RECT  1.450 1.600 1.690 2.360 ;
        RECT  1.450 2.120 3.240 2.360 ;
        RECT  3.000 2.120 3.240 2.770 ;
        RECT  2.000 2.120 2.240 3.460 ;
        RECT  0.930 3.220 2.240 3.460 ;
        RECT  2.730 1.640 3.960 1.880 ;
        RECT  3.550 1.640 3.960 2.080 ;
        RECT  2.480 3.220 3.790 3.460 ;
        RECT  3.550 1.640 3.790 3.600 ;
        RECT  3.390 3.220 3.790 3.600 ;
        RECT  4.000 1.060 4.470 1.380 ;
        RECT  4.200 1.060 4.470 3.440 ;
        RECT  4.030 3.200 4.300 4.130 ;
        RECT  5.520 1.150 5.800 1.710 ;
        RECT  5.520 1.150 5.760 4.130 ;
        RECT  6.000 3.280 6.860 3.520 ;
        RECT  4.820 1.150 5.060 4.610 ;
        RECT  4.780 3.640 5.060 4.610 ;
        RECT  6.000 3.280 6.240 4.610 ;
        RECT  4.780 4.370 6.240 4.610 ;
        RECT  7.040 1.300 7.340 2.150 ;
        RECT  6.000 1.910 7.340 2.150 ;
        RECT  7.100 1.300 7.340 4.130 ;
        RECT  6.800 3.810 7.340 4.130 ;
    END
END lanhn2

MACRO lanhn1
    CLASS CORE ;
    FOREIGN lanhn1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.700 2.740 4.200 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.480 ;
        END
    END E
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.500  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.380 1.110 8.840 2.490 ;
        RECT  8.380 1.110 8.620 3.450 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.610 4.130 7.850 5.600 ;
        RECT  6.470 4.710 6.870 5.600 ;
        RECT  3.300 3.840 3.540 5.600 ;
        RECT  1.780 3.700 2.020 5.600 ;
        RECT  0.420 4.710 0.820 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.500 0.000 7.900 0.980 ;
        RECT  6.320 0.000 6.560 1.550 ;
        RECT  3.330 0.000 3.570 1.200 ;
        RECT  2.220 0.000 2.460 1.200 ;
        RECT  0.720 0.000 0.960 1.210 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 2.600 1.760 2.840 ;
        RECT  0.740 1.550 0.980 2.960 ;
        RECT  0.440 2.720 0.980 2.960 ;
        RECT  0.440 2.720 0.680 4.370 ;
        RECT  0.440 4.050 0.820 4.370 ;
        RECT  1.450 1.600 1.690 2.360 ;
        RECT  1.450 2.120 3.240 2.360 ;
        RECT  3.000 2.120 3.240 2.770 ;
        RECT  2.000 2.120 2.240 3.460 ;
        RECT  0.930 3.220 2.240 3.460 ;
        RECT  2.730 1.640 3.980 1.880 ;
        RECT  3.550 1.640 3.980 2.080 ;
        RECT  2.480 3.220 3.790 3.460 ;
        RECT  3.550 1.640 3.790 3.600 ;
        RECT  3.390 3.220 3.790 3.600 ;
        RECT  4.020 1.060 4.490 1.380 ;
        RECT  4.220 1.060 4.490 3.440 ;
        RECT  4.030 3.200 4.300 4.130 ;
        RECT  5.580 1.150 5.820 3.040 ;
        RECT  5.520 2.800 5.760 4.130 ;
        RECT  6.000 3.280 6.860 3.520 ;
        RECT  4.840 1.150 5.080 4.610 ;
        RECT  4.780 3.640 5.080 4.610 ;
        RECT  6.000 3.280 6.240 4.610 ;
        RECT  4.780 4.370 6.240 4.610 ;
        RECT  7.070 1.300 7.340 2.150 ;
        RECT  6.060 1.910 7.340 2.150 ;
        RECT  7.100 1.300 7.340 4.130 ;
        RECT  6.800 3.810 7.340 4.130 ;
    END
END lanhn1

MACRO lanhb4
    CLASS CORE ;
    FOREIGN lanhb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.260 2.290 2.740 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.380  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.260 0.700 3.020 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.346  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.060 1.690 10.580 2.710 ;
        RECT  8.860 4.020 10.480 4.340 ;
        RECT  10.060 1.690 10.480 4.340 ;
        RECT  9.980 1.690 10.580 2.090 ;
        RECT  8.860 3.660 9.100 4.340 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.515  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.120 1.120 8.520 1.520 ;
        RECT  8.060 1.220 8.460 2.460 ;
        RECT  6.260 3.330 8.070 3.730 ;
        RECT  7.650 2.020 8.070 3.730 ;
        RECT  7.120 1.220 8.520 1.460 ;
        RECT  6.640 1.200 7.270 1.440 ;
        RECT  6.260 3.010 6.500 3.730 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  10.720 3.260 10.960 5.600 ;
        RECT  9.340 4.590 9.740 5.600 ;
        RECT  8.040 4.590 8.440 5.600 ;
        RECT  6.570 4.620 6.970 5.600 ;
        RECT  4.730 4.340 5.130 5.600 ;
        RECT  2.160 4.540 2.560 5.600 ;
        RECT  0.750 4.230 1.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  10.540 0.000 10.940 1.150 ;
        RECT  8.860 0.000 9.260 0.980 ;
        RECT  7.380 0.000 7.780 0.980 ;
        RECT  5.200 0.000 5.600 1.420 ;
        RECT  2.210 1.580 2.780 1.820 ;
        RECT  2.540 0.000 2.780 1.820 ;
        RECT  0.490 0.000 0.890 0.930 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.760 1.180 2.000 ;
        RECT  0.940 2.490 1.480 2.890 ;
        RECT  0.940 1.760 1.180 3.580 ;
        RECT  0.150 3.340 1.180 3.580 ;
        RECT  1.540 0.980 2.100 1.220 ;
        RECT  1.540 0.980 1.780 1.650 ;
        RECT  1.590 1.500 1.830 2.260 ;
        RECT  1.780 2.020 2.020 4.010 ;
        RECT  1.450 3.610 2.020 4.010 ;
        RECT  3.030 1.500 3.270 2.260 ;
        RECT  2.980 2.010 3.220 4.120 ;
        RECT  2.750 3.720 3.220 4.120 ;
        RECT  4.280 1.200 4.860 1.440 ;
        RECT  4.280 1.200 4.520 3.570 ;
        RECT  4.120 3.170 4.520 3.570 ;
        RECT  6.020 1.120 6.260 2.060 ;
        RECT  6.020 1.710 7.280 2.060 ;
        RECT  4.760 1.820 7.280 2.060 ;
        RECT  6.340 1.710 7.280 2.110 ;
        RECT  4.760 1.820 5.160 2.220 ;
        RECT  5.770 1.820 6.010 3.560 ;
        RECT  5.470 3.160 6.010 3.560 ;
        RECT  3.800 1.290 4.040 2.680 ;
        RECT  3.460 2.440 4.040 2.680 ;
        RECT  5.130 2.500 5.530 2.900 ;
        RECT  8.700 2.520 9.650 2.920 ;
        RECT  8.380 2.700 8.890 3.010 ;
        RECT  3.460 2.440 3.700 4.100 ;
        RECT  4.990 2.680 5.230 4.100 ;
        RECT  3.460 3.860 5.900 4.100 ;
        RECT  8.380 2.700 8.620 4.290 ;
        RECT  5.650 4.050 8.620 4.290 ;
    END
END lanhb4

MACRO lanhb2
    CLASS CORE ;
    FOREIGN lanhb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.990 3.580 ;
        RECT  2.710 2.030 2.990 3.580 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.450 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.322  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.150 3.050 7.780 3.580 ;
        RECT  7.420 1.380 7.660 3.580 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.322  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.460 3.050 9.080 3.580 ;
        RECT  8.840 1.380 9.080 3.580 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  9.450 4.060 9.690 5.600 ;
        RECT  7.970 4.060 8.210 5.600 ;
        RECT  6.490 4.060 6.730 5.600 ;
        RECT  5.160 4.170 5.400 5.600 ;
        RECT  2.290 4.400 2.530 5.600 ;
        RECT  0.630 4.510 1.030 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  9.450 0.000 9.850 0.890 ;
        RECT  8.060 0.000 8.460 0.890 ;
        RECT  6.670 0.000 7.070 0.890 ;
        RECT  5.250 0.000 5.650 0.890 ;
        RECT  2.200 0.000 2.600 0.890 ;
        RECT  0.670 0.000 1.070 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.780 1.460 1.380 1.700 ;
        RECT  1.140 1.460 1.380 4.090 ;
        RECT  0.810 3.850 1.380 4.090 ;
        RECT  1.660 2.470 2.140 2.870 ;
        RECT  1.660 1.500 1.900 4.080 ;
        RECT  2.950 1.540 3.510 1.780 ;
        RECT  3.270 1.540 3.510 4.060 ;
        RECT  2.930 3.820 3.510 4.060 ;
        RECT  4.560 1.500 4.800 3.450 ;
        RECT  5.040 2.600 6.170 2.840 ;
        RECT  3.820 1.500 4.060 4.270 ;
        RECT  5.040 2.600 5.280 3.930 ;
        RECT  3.820 3.690 5.280 3.930 ;
        RECT  3.820 3.690 4.090 4.270 ;
        RECT  6.100 1.500 6.340 2.350 ;
        RECT  5.040 2.110 6.650 2.350 ;
        RECT  6.410 2.110 6.650 3.370 ;
        RECT  5.820 3.130 6.650 3.370 ;
    END
END lanhb2

MACRO lanhb1
    CLASS CORE ;
    FOREIGN lanhb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 3.070 3.580 ;
        RECT  2.830 2.020 3.070 3.580 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.247  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.450 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.141  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.010 2.020 7.780 2.460 ;
        RECT  7.010 1.460 7.250 4.130 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.165  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.430 1.460 8.840 3.450 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.750 4.060 7.990 5.600 ;
        RECT  5.640 4.240 5.880 5.600 ;
        RECT  2.360 4.390 2.600 5.600 ;
        RECT  0.630 4.510 1.030 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.670 0.000 8.070 0.890 ;
        RECT  5.390 0.000 5.790 0.890 ;
        RECT  2.350 0.000 2.750 0.890 ;
        RECT  0.670 0.000 1.070 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.780 1.460 1.380 1.700 ;
        RECT  1.140 1.460 1.380 4.090 ;
        RECT  0.810 3.850 1.380 4.090 ;
        RECT  1.700 1.500 2.020 2.870 ;
        RECT  1.700 2.470 2.140 2.870 ;
        RECT  1.700 1.500 1.940 4.100 ;
        RECT  3.080 1.540 3.710 1.780 ;
        RECT  3.470 1.540 3.710 4.100 ;
        RECT  3.090 3.860 3.710 4.100 ;
        RECT  4.690 1.500 4.930 3.520 ;
        RECT  4.690 3.200 5.190 3.520 ;
        RECT  3.950 1.500 4.190 4.480 ;
        RECT  5.890 2.590 6.130 4.000 ;
        RECT  3.950 3.760 6.130 4.000 ;
        RECT  3.950 3.760 4.210 4.480 ;
        RECT  6.240 1.500 6.480 2.350 ;
        RECT  5.170 2.110 6.620 2.350 ;
        RECT  6.380 2.110 6.620 3.520 ;
    END
END lanhb1

MACRO laclq4
    CLASS CORE ;
    FOREIGN laclq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.979  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 1.460 6.100 1.900 ;
        RECT  5.660 0.980 5.900 2.530 ;
        RECT  2.720 0.980 5.900 1.220 ;
        RECT  3.180 2.040 3.420 2.920 ;
        RECT  2.720 2.040 3.420 2.280 ;
        RECT  2.720 0.980 2.960 2.280 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.451  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.520 2.800 3.020 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.800 2.840 ;
        RECT  0.120 2.580 0.500 3.020 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.050  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.560 3.320 10.580 3.560 ;
        RECT  10.340 1.690 10.580 3.560 ;
        RECT  10.140 2.580 10.580 3.020 ;
        RECT  8.420 1.690 10.580 1.930 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  10.530 4.620 10.930 5.600 ;
        RECT  9.120 4.610 9.520 5.600 ;
        RECT  7.820 4.610 8.220 5.600 ;
        RECT  5.750 4.270 5.990 5.600 ;
        RECT  2.800 4.710 3.200 5.600 ;
        RECT  0.880 4.290 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  9.190 0.000 9.590 0.890 ;
        RECT  7.650 0.000 8.050 0.890 ;
        RECT  6.390 0.000 6.790 0.890 ;
        RECT  2.030 0.000 2.430 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.580 1.350 1.820 ;
        RECT  1.110 1.580 1.350 2.260 ;
        RECT  1.180 2.020 1.420 2.860 ;
        RECT  1.040 2.620 1.280 3.500 ;
        RECT  0.150 3.260 1.280 3.500 ;
        RECT  3.260 1.480 3.900 1.720 ;
        RECT  3.660 1.480 3.900 3.660 ;
        RECT  2.150 3.420 3.900 3.660 ;
        RECT  2.150 3.420 2.550 3.820 ;
        RECT  1.590 1.230 1.830 1.780 ;
        RECT  1.660 1.540 1.900 3.340 ;
        RECT  1.530 3.100 1.770 4.300 ;
        RECT  2.810 3.900 4.380 4.140 ;
        RECT  4.140 2.520 4.380 4.140 ;
        RECT  1.530 4.060 3.050 4.300 ;
        RECT  4.800 1.460 5.420 1.700 ;
        RECT  5.180 2.820 6.770 3.060 ;
        RECT  5.180 1.460 5.420 3.450 ;
        RECT  6.530 2.820 6.770 3.480 ;
        RECT  7.050 1.650 7.430 2.050 ;
        RECT  6.280 2.310 7.430 2.550 ;
        RECT  7.190 1.650 7.430 3.450 ;
        RECT  7.190 3.050 7.650 3.450 ;
        RECT  4.140 1.460 4.380 2.280 ;
        RECT  4.140 2.040 4.860 2.280 ;
        RECT  7.670 2.410 9.690 2.810 ;
        RECT  7.890 2.410 8.130 4.030 ;
        RECT  4.620 3.790 8.130 4.030 ;
        RECT  4.620 2.040 4.860 4.620 ;
        RECT  4.190 4.380 4.860 4.620 ;
    END
END laclq4

MACRO laclq2
    CLASS CORE ;
    FOREIGN laclq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.020 1.370 2.480 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.340  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.830 0.500 3.580 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.207  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.470 3.020 ;
        RECT  2.230 2.090 2.470 3.020 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.790 1.460 9.460 1.900 ;
        RECT  8.790 1.140 9.190 1.900 ;
        RECT  8.790 1.140 9.080 3.550 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  9.530 4.710 9.930 5.600 ;
        RECT  7.980 4.710 8.380 5.600 ;
        RECT  6.030 4.710 6.430 5.600 ;
        RECT  2.560 4.710 2.960 5.600 ;
        RECT  1.510 4.710 1.910 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  9.530 0.000 9.930 1.010 ;
        RECT  8.040 0.000 8.440 1.010 ;
        RECT  6.830 0.000 7.070 1.540 ;
        RECT  2.680 0.000 3.080 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.910 1.610 3.030 1.850 ;
        RECT  2.790 2.090 3.310 2.480 ;
        RECT  2.790 1.610 3.030 3.500 ;
        RECT  1.970 3.260 3.030 3.500 ;
        RECT  3.270 1.610 3.910 1.850 ;
        RECT  3.670 1.610 3.910 3.460 ;
        RECT  3.330 3.220 3.910 3.460 ;
        RECT  3.970 1.050 4.400 1.370 ;
        RECT  1.200 1.130 4.400 1.370 ;
        RECT  1.200 1.130 1.520 1.630 ;
        RECT  0.740 3.750 1.060 4.260 ;
        RECT  4.160 1.050 4.400 4.260 ;
        RECT  0.740 4.020 4.400 4.260 ;
        RECT  5.530 1.440 5.770 3.780 ;
        RECT  5.340 3.460 7.120 3.780 ;
        RECT  6.500 2.050 7.770 2.290 ;
        RECT  7.530 1.720 7.770 3.550 ;
        RECT  7.500 2.050 7.770 3.550 ;
        RECT  4.690 1.440 5.110 1.760 ;
        RECT  4.690 1.440 4.930 4.260 ;
        RECT  8.060 2.620 8.300 4.260 ;
        RECT  4.690 4.020 8.300 4.260 ;
    END
END laclq2

MACRO laclq1
    CLASS CORE ;
    FOREIGN laclq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.344  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 1.420 2.940 ;
        RECT  0.620 2.020 1.420 2.460 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.700 0.800 3.020 ;
        RECT  0.120 2.700 0.500 3.580 ;
        END
    END D
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.230 2.630 2.470 ;
        RECT  1.740 2.230 2.180 3.020 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.264  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.050 1.710 9.400 3.620 ;
        RECT  8.900 1.710 9.400 2.460 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  8.200 4.710 8.600 5.600 ;
        RECT  6.240 4.710 6.640 5.600 ;
        RECT  2.660 4.710 3.060 5.600 ;
        RECT  1.570 4.710 1.970 5.600 ;
        RECT  0.170 4.710 0.570 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.210 0.000 8.450 1.370 ;
        RECT  6.920 0.000 7.160 1.490 ;
        RECT  2.870 0.000 3.270 0.890 ;
        RECT  0.230 0.000 0.470 1.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.070 1.610 3.110 1.850 ;
        RECT  2.870 2.220 3.430 2.460 ;
        RECT  2.870 1.610 3.110 3.500 ;
        RECT  2.070 3.260 3.110 3.500 ;
        RECT  3.460 1.610 4.000 1.930 ;
        RECT  3.760 1.610 4.000 2.970 ;
        RECT  3.760 2.570 4.110 2.970 ;
        RECT  3.510 2.730 4.110 2.970 ;
        RECT  3.510 2.730 3.750 3.540 ;
        RECT  4.160 1.050 4.590 1.370 ;
        RECT  1.350 1.130 4.590 1.370 ;
        RECT  1.350 1.130 1.750 1.530 ;
        RECT  4.130 3.220 4.590 4.020 ;
        RECT  4.350 1.050 4.590 4.020 ;
        RECT  0.800 3.780 4.590 4.020 ;
        RECT  5.720 1.230 5.960 3.620 ;
        RECT  5.610 3.300 7.330 3.540 ;
        RECT  5.610 3.300 6.010 3.620 ;
        RECT  7.540 1.770 7.950 2.270 ;
        RECT  6.590 2.030 7.950 2.270 ;
        RECT  7.710 1.770 7.950 3.620 ;
        RECT  4.950 1.230 5.310 1.630 ;
        RECT  4.950 1.230 5.190 4.100 ;
        RECT  8.290 2.690 8.530 4.100 ;
        RECT  4.950 3.860 8.530 4.100 ;
    END
END laclq1

MACRO lachq4
    CLASS CORE ;
    FOREIGN lachq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.504  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.110 2.020 6.660 2.460 ;
        RECT  6.110 2.020 6.350 2.860 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.260 2.580 2.970 3.020 ;
        RECT  2.730 2.260 2.970 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 1.900 ;
        RECT  0.600 2.310 1.420 2.550 ;
        RECT  1.180 1.460 1.420 2.550 ;
        RECT  0.600 2.310 0.840 2.950 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.060  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.500 3.020 11.080 3.260 ;
        RECT  10.620 1.360 11.080 3.260 ;
        RECT  8.880 1.360 11.080 1.770 ;
        RECT  9.800 3.020 10.040 4.180 ;
        RECT  8.500 3.020 8.740 4.580 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  10.460 4.300 10.860 5.600 ;
        RECT  9.060 3.500 9.300 5.600 ;
        RECT  7.620 4.180 8.020 5.600 ;
        RECT  5.660 4.700 6.060 5.600 ;
        RECT  2.910 4.700 3.310 5.600 ;
        RECT  0.800 4.700 1.200 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  9.680 0.000 10.080 1.120 ;
        RECT  8.150 0.000 8.550 1.370 ;
        RECT  6.530 1.010 7.100 1.250 ;
        RECT  6.860 0.000 7.100 1.250 ;
        RECT  2.160 0.000 2.560 0.890 ;
        RECT  0.920 0.000 1.320 0.900 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.140 0.980 0.690 1.220 ;
        RECT  0.450 0.980 0.690 2.070 ;
        RECT  0.120 1.660 0.690 2.070 ;
        RECT  0.120 1.660 0.360 3.730 ;
        RECT  1.280 2.790 1.520 3.640 ;
        RECT  0.120 3.400 1.520 3.640 ;
        RECT  0.120 3.320 0.590 3.730 ;
        RECT  3.350 1.460 3.910 1.700 ;
        RECT  3.350 1.460 3.590 3.460 ;
        RECT  3.180 3.220 3.900 3.460 ;
        RECT  2.340 3.420 2.580 3.970 ;
        RECT  3.180 3.220 3.420 3.970 ;
        RECT  2.340 3.730 3.420 3.970 ;
        RECT  3.660 3.220 3.900 3.970 ;
        RECT  2.870 0.980 4.390 1.220 ;
        RECT  1.860 1.150 3.110 1.390 ;
        RECT  4.150 0.980 4.390 2.300 ;
        RECT  3.920 1.960 4.390 2.300 ;
        RECT  1.860 1.150 2.100 2.340 ;
        RECT  1.760 2.100 2.000 3.620 ;
        RECT  5.150 2.330 5.390 3.680 ;
        RECT  4.290 3.440 5.390 3.680 ;
        RECT  1.850 2.100 2.000 4.120 ;
        RECT  1.490 3.880 2.100 4.120 ;
        RECT  1.860 3.390 2.100 4.460 ;
        RECT  4.290 3.440 4.540 4.460 ;
        RECT  1.860 4.210 4.540 4.460 ;
        RECT  5.400 1.840 5.790 2.090 ;
        RECT  5.400 1.500 5.640 2.090 ;
        RECT  5.550 1.910 5.870 2.150 ;
        RECT  5.630 1.910 5.870 4.190 ;
        RECT  4.950 3.950 6.740 4.190 ;
        RECT  4.630 1.020 6.270 1.260 ;
        RECT  6.030 1.490 6.480 1.730 ;
        RECT  6.030 1.020 6.270 1.730 ;
        RECT  6.240 1.540 7.140 1.780 ;
        RECT  6.900 1.540 7.140 2.440 ;
        RECT  6.900 2.200 7.820 2.440 ;
        RECT  4.630 1.020 4.870 3.200 ;
        RECT  4.200 2.960 4.870 3.200 ;
        RECT  7.470 1.280 7.710 1.960 ;
        RECT  7.470 1.720 8.300 1.960 ;
        RECT  8.060 1.720 8.300 2.880 ;
        RECT  6.720 2.700 8.270 2.940 ;
        RECT  7.080 2.700 7.530 3.540 ;
    END
END lachq4

MACRO lachq2
    CLASS CORE ;
    FOREIGN lachq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.220 2.090 1.620 3.580 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.496  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.490 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.160 2.740 3.020 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.277  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.850 2.020 9.460 2.460 ;
        RECT  8.850 1.460 9.170 2.460 ;
        RECT  8.850 1.460 9.090 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  9.580 4.060 9.820 5.600 ;
        RECT  8.140 4.710 8.540 5.600 ;
        RECT  6.080 4.710 6.480 5.600 ;
        RECT  2.760 4.550 3.160 5.600 ;
        RECT  1.460 4.550 1.860 5.600 ;
        RECT  0.150 4.550 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  9.610 0.000 9.850 1.300 ;
        RECT  8.160 0.000 8.560 1.080 ;
        RECT  6.900 0.000 7.300 1.110 ;
        RECT  2.930 0.000 3.170 1.360 ;
        RECT  0.210 0.000 0.610 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.110 1.680 3.220 1.920 ;
        RECT  2.980 2.820 3.340 3.220 ;
        RECT  2.980 1.680 3.220 3.750 ;
        RECT  1.990 3.510 3.220 3.750 ;
        RECT  3.460 1.630 3.820 1.950 ;
        RECT  3.580 2.430 4.080 2.830 ;
        RECT  3.580 1.630 3.820 3.830 ;
        RECT  3.460 3.430 3.820 3.830 ;
        RECT  0.740 1.610 1.810 1.850 ;
        RECT  4.170 1.850 4.720 2.090 ;
        RECT  0.740 1.610 0.980 2.970 ;
        RECT  4.480 1.850 4.720 3.310 ;
        RECT  4.210 3.070 4.720 3.310 ;
        RECT  0.700 2.730 0.940 4.310 ;
        RECT  0.700 3.830 1.120 4.310 ;
        RECT  0.700 4.070 4.450 4.310 ;
        RECT  4.210 3.070 4.450 4.600 ;
        RECT  3.990 4.070 4.450 4.600 ;
        RECT  5.730 1.770 5.970 3.060 ;
        RECT  5.550 2.820 5.790 3.990 ;
        RECT  5.550 3.750 7.250 3.990 ;
        RECT  7.500 1.460 7.750 2.620 ;
        RECT  6.600 2.380 7.790 2.620 ;
        RECT  7.550 2.380 7.790 3.450 ;
        RECT  4.990 1.770 5.230 3.790 ;
        RECT  4.810 3.550 5.050 4.470 ;
        RECT  8.300 2.520 8.540 4.470 ;
        RECT  4.810 4.230 8.540 4.470 ;
    END
END lachq2

MACRO lachq1
    CLASS CORE ;
    FOREIGN lachq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.220 2.090 1.620 3.580 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.496  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.490 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.100 2.740 3.020 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.000  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 1.460 9.400 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  8.370 4.710 8.770 5.600 ;
        RECT  6.240 4.710 6.640 5.600 ;
        RECT  2.760 4.550 3.160 5.600 ;
        RECT  1.460 4.550 1.860 5.600 ;
        RECT  0.150 4.550 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.320 0.000 8.720 1.080 ;
        RECT  6.960 0.000 7.200 1.710 ;
        RECT  2.930 0.000 3.170 1.370 ;
        RECT  0.210 0.000 0.610 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.190 1.000 2.430 1.850 ;
        RECT  2.190 1.610 3.220 1.850 ;
        RECT  2.980 2.670 3.440 3.070 ;
        RECT  2.980 1.610 3.220 3.750 ;
        RECT  2.110 3.510 3.220 3.750 ;
        RECT  3.460 1.630 3.930 1.950 ;
        RECT  3.660 1.630 3.930 2.570 ;
        RECT  3.730 2.430 4.180 2.830 ;
        RECT  3.730 2.430 3.980 3.830 ;
        RECT  3.570 3.430 3.980 3.830 ;
        RECT  0.740 1.380 1.810 1.620 ;
        RECT  4.170 1.770 4.660 2.090 ;
        RECT  0.740 1.380 0.980 2.970 ;
        RECT  0.700 2.730 0.940 4.310 ;
        RECT  0.700 3.830 1.120 4.310 ;
        RECT  0.700 4.070 4.660 4.310 ;
        RECT  4.420 1.770 4.660 4.600 ;
        RECT  4.150 4.070 4.660 4.600 ;
        RECT  5.710 1.770 5.970 3.990 ;
        RECT  5.710 3.750 7.410 3.990 ;
        RECT  7.660 1.460 7.900 2.620 ;
        RECT  6.760 2.380 7.950 2.620 ;
        RECT  7.710 2.380 7.950 3.450 ;
        RECT  4.970 1.770 5.230 4.470 ;
        RECT  8.300 2.520 8.540 4.470 ;
        RECT  4.970 4.230 8.540 4.470 ;
    END
END lachq1

MACRO labhb4
    CLASS CORE ;
    FOREIGN labhb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.250 2.570 3.860 3.020 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.433  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.150 2.550 2.740 3.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.451  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.600 0.930 3.000 ;
        RECT  0.120 1.880 0.500 3.000 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.981  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.590 3.360 12.310 3.600 ;
        RECT  10.400 1.240 12.280 1.480 ;
        RECT  11.260 3.140 11.700 3.600 ;
        RECT  11.420 1.240 11.660 3.600 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.700  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.510 2.780 14.910 3.320 ;
        RECT  14.060 1.460 14.600 1.900 ;
        RECT  13.370 2.780 14.910 3.020 ;
        RECT  13.040 1.570 14.600 1.810 ;
        RECT  13.210 3.940 13.610 4.350 ;
        RECT  13.370 1.570 13.610 4.350 ;
        RECT  13.040 0.980 13.280 1.810 ;
        RECT  12.710 0.980 13.280 1.220 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.506  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.440 2.020 8.900 2.460 ;
        RECT  8.440 2.020 8.680 2.840 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  15.200 3.550 15.470 5.600 ;
        RECT  13.850 3.260 14.090 5.600 ;
        RECT  12.650 4.620 13.050 5.600 ;
        RECT  11.350 4.320 11.750 5.600 ;
        RECT  10.050 4.320 10.450 5.600 ;
        RECT  7.870 4.290 8.270 5.600 ;
        RECT  6.030 4.370 6.430 5.600 ;
        RECT  2.730 4.330 3.130 5.600 ;
        RECT  0.720 4.400 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  15.020 0.000 15.260 1.780 ;
        RECT  13.540 0.000 13.780 1.330 ;
        RECT  11.140 0.000 11.540 0.980 ;
        RECT  9.740 0.000 9.980 1.370 ;
        RECT  8.370 0.000 8.770 0.890 ;
        RECT  6.510 0.000 6.910 0.890 ;
        RECT  2.270 0.000 2.670 1.010 ;
        RECT  0.720 0.000 1.120 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.130 1.760 1.370 ;
        RECT  1.360 0.980 1.760 1.380 ;
        RECT  0.230 1.130 0.630 1.640 ;
        RECT  1.190 1.130 1.430 3.490 ;
        RECT  0.150 3.250 1.430 3.490 ;
        RECT  3.440 1.690 3.680 2.330 ;
        RECT  3.440 2.090 4.340 2.330 ;
        RECT  4.100 2.090 4.340 3.500 ;
        RECT  2.160 3.260 4.340 3.500 ;
        RECT  2.960 0.980 4.010 1.220 ;
        RECT  2.960 0.980 3.200 1.860 ;
        RECT  1.670 1.620 3.200 1.860 ;
        RECT  1.670 3.850 3.610 4.090 ;
        RECT  5.060 2.740 5.300 4.140 ;
        RECT  3.370 3.900 5.300 4.140 ;
        RECT  1.670 1.620 1.910 4.620 ;
        RECT  1.460 4.220 1.910 4.620 ;
        RECT  4.580 1.140 7.910 1.380 ;
        RECT  4.100 1.610 4.820 1.850 ;
        RECT  7.670 1.140 7.910 2.670 ;
        RECT  7.320 2.430 7.910 2.670 ;
        RECT  4.580 1.140 4.820 3.660 ;
        RECT  6.300 1.620 7.430 1.860 ;
        RECT  6.300 1.620 6.540 3.210 ;
        RECT  6.300 2.970 7.550 3.210 ;
        RECT  7.300 3.140 9.010 3.380 ;
        RECT  7.300 3.120 7.700 3.530 ;
        RECT  9.000 1.540 9.380 1.780 ;
        RECT  9.000 1.160 9.240 1.780 ;
        RECT  9.140 1.770 11.180 2.010 ;
        RECT  9.390 1.770 9.630 3.470 ;
        RECT  5.060 1.620 5.300 2.290 ;
        RECT  5.060 2.050 5.780 2.290 ;
        RECT  6.680 3.450 6.920 4.130 ;
        RECT  6.680 3.810 8.900 4.050 ;
        RECT  12.550 1.710 12.790 4.080 ;
        RECT  8.510 3.840 12.790 4.080 ;
        RECT  5.540 3.890 6.930 4.130 ;
        RECT  5.540 2.050 5.780 4.620 ;
        RECT  5.220 4.380 5.780 4.620 ;
        RECT  13.910 2.140 16.010 2.540 ;
        RECT  15.770 1.480 16.010 4.620 ;
    END
END labhb4

MACRO labhb2
    CLASS CORE ;
    FOREIGN labhb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.100 1.500 3.580 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.800 2.840 ;
        RECT  0.120 2.020 0.500 2.840 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.207  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.020 2.810 2.460 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.322  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.380 3.140 12.950 3.580 ;
        RECT  12.380 1.380 12.740 3.580 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.322  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.070 3.130 11.700 3.580 ;
        RECT  11.070 1.380 11.320 3.580 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.360  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.580 7.670 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.120 5.600 ;
        RECT  14.280 4.170 14.520 5.600 ;
        RECT  13.370 4.060 13.610 5.600 ;
        RECT  11.890 4.060 12.130 5.600 ;
        RECT  10.410 4.130 10.650 5.600 ;
        RECT  9.280 4.200 9.520 5.600 ;
        RECT  7.800 4.220 8.040 5.600 ;
        RECT  6.420 4.220 6.660 5.600 ;
        RECT  2.830 4.220 3.070 5.600 ;
        RECT  1.740 4.300 1.980 5.600 ;
        RECT  0.230 4.220 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.120 0.740 ;
        RECT  14.150 0.000 14.550 1.060 ;
        RECT  13.190 0.000 13.430 1.230 ;
        RECT  11.800 0.000 12.040 1.230 ;
        RECT  10.330 0.000 10.730 1.050 ;
        RECT  9.550 0.000 9.950 1.080 ;
        RECT  6.950 0.000 7.350 1.130 ;
        RECT  2.760 0.000 3.160 1.040 ;
        RECT  1.730 0.000 2.150 0.820 ;
        RECT  0.230 0.000 0.470 1.600 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.170 1.460 3.290 1.700 ;
        RECT  3.050 1.460 3.290 2.940 ;
        RECT  3.050 2.530 3.510 2.940 ;
        RECT  2.240 2.700 3.510 2.940 ;
        RECT  2.240 2.700 2.480 3.500 ;
        RECT  3.530 1.460 3.990 1.860 ;
        RECT  3.750 2.030 4.190 2.430 ;
        RECT  3.750 1.460 3.990 3.500 ;
        RECT  3.520 3.180 3.990 3.500 ;
        RECT  4.230 1.390 4.680 1.790 ;
        RECT  1.430 1.450 1.670 2.580 ;
        RECT  1.430 2.340 1.980 2.580 ;
        RECT  4.440 1.390 4.680 3.080 ;
        RECT  4.300 2.840 4.540 3.980 ;
        RECT  1.740 3.740 4.540 3.980 ;
        RECT  1.740 2.340 1.980 4.060 ;
        RECT  0.890 3.820 1.980 4.060 ;
        RECT  7.680 1.070 9.020 1.310 ;
        RECT  7.680 1.070 7.920 1.610 ;
        RECT  5.690 1.370 7.920 1.610 ;
        RECT  5.690 1.370 6.030 3.500 ;
        RECT  5.690 3.260 7.420 3.500 ;
        RECT  7.940 3.190 9.050 3.430 ;
        RECT  5.040 1.370 5.290 3.980 ;
        RECT  7.940 3.190 8.180 3.980 ;
        RECT  5.040 3.740 8.180 3.980 ;
        RECT  7.240 1.850 9.000 2.090 ;
        RECT  6.650 1.980 7.480 2.220 ;
        RECT  8.760 1.850 9.000 2.950 ;
        RECT  8.760 2.710 9.530 2.950 ;
        RECT  9.290 2.710 9.530 3.960 ;
        RECT  8.460 3.720 9.530 3.960 ;
        RECT  9.290 1.430 9.530 2.450 ;
        RECT  9.290 2.210 10.410 2.450 ;
        RECT  9.880 2.210 10.410 2.610 ;
        RECT  9.880 2.210 10.120 3.710 ;
        RECT  12.980 2.290 14.430 2.530 ;
        RECT  14.190 1.410 14.430 3.830 ;
    END
END labhb2

MACRO labhb1
    CLASS CORE ;
    FOREIGN labhb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.100 1.500 3.580 ;
        END
    END CDN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.530 0.800 2.850 ;
        RECT  0.120 2.020 0.500 2.850 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.207  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.020 2.810 2.460 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.085  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.200 3.130 12.370 3.370 ;
        RECT  11.200 1.460 12.330 1.900 ;
        RECT  11.200 1.460 11.440 3.370 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.650 1.460 10.890 3.450 ;
        RECT  10.140 1.460 10.890 1.940 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.360  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.580 7.670 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 14.000 5.600 ;
        RECT  12.940 4.170 13.180 5.600 ;
        RECT  11.390 4.080 11.630 5.600 ;
        RECT  9.280 4.200 9.520 5.600 ;
        RECT  7.800 4.220 8.040 5.600 ;
        RECT  6.420 4.220 6.660 5.600 ;
        RECT  2.830 4.220 3.070 5.600 ;
        RECT  1.740 4.300 1.980 5.600 ;
        RECT  0.230 4.220 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 14.000 0.740 ;
        RECT  12.980 0.000 13.380 1.060 ;
        RECT  11.160 0.000 11.560 1.220 ;
        RECT  9.660 0.000 10.060 1.080 ;
        RECT  6.950 0.000 7.350 1.130 ;
        RECT  2.760 0.000 3.160 0.890 ;
        RECT  1.730 0.000 2.150 0.820 ;
        RECT  0.230 0.000 0.470 1.600 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.170 1.460 3.290 1.700 ;
        RECT  3.050 1.460 3.290 2.940 ;
        RECT  3.050 2.530 3.510 2.940 ;
        RECT  2.240 2.700 3.510 2.940 ;
        RECT  2.240 2.700 2.480 3.500 ;
        RECT  3.530 1.460 3.990 1.860 ;
        RECT  3.750 2.030 4.190 2.430 ;
        RECT  3.750 1.460 3.990 3.500 ;
        RECT  3.520 3.180 3.990 3.500 ;
        RECT  4.230 1.390 4.680 1.790 ;
        RECT  1.430 1.450 1.670 2.580 ;
        RECT  1.430 2.340 1.980 2.580 ;
        RECT  4.440 1.390 4.680 3.080 ;
        RECT  4.300 2.840 4.540 3.980 ;
        RECT  1.740 3.740 4.540 3.980 ;
        RECT  1.740 2.340 1.980 4.060 ;
        RECT  0.890 3.820 1.980 4.060 ;
        RECT  7.680 1.070 9.020 1.310 ;
        RECT  7.680 1.070 7.920 1.610 ;
        RECT  5.690 1.370 7.920 1.610 ;
        RECT  5.690 1.370 6.030 3.500 ;
        RECT  5.690 3.260 7.420 3.500 ;
        RECT  7.940 3.190 9.050 3.430 ;
        RECT  5.040 1.370 5.290 3.980 ;
        RECT  7.940 3.190 8.180 3.980 ;
        RECT  5.040 3.740 8.180 3.980 ;
        RECT  7.240 1.850 9.000 2.090 ;
        RECT  6.650 1.980 7.480 2.220 ;
        RECT  8.760 1.850 9.000 2.950 ;
        RECT  8.760 2.710 9.530 2.950 ;
        RECT  9.290 2.710 9.530 3.960 ;
        RECT  8.460 3.720 9.530 3.960 ;
        RECT  9.400 1.430 9.640 2.450 ;
        RECT  9.400 2.210 10.410 2.450 ;
        RECT  9.880 2.210 10.410 2.610 ;
        RECT  9.880 2.210 10.120 3.710 ;
        RECT  11.680 2.150 13.090 2.390 ;
        RECT  12.850 1.410 13.090 3.830 ;
    END
END labhb1

MACRO jkbrb4
    CLASS CORE ;
    FOREIGN jkbrb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.710  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.470 1.130 15.710 2.520 ;
        RECT  13.390 1.130 15.710 1.370 ;
        RECT  9.790 0.980 13.620 1.220 ;
        RECT  9.210 1.500 10.030 1.740 ;
        RECT  9.790 0.980 10.030 1.740 ;
        RECT  9.020 2.020 9.460 2.460 ;
        RECT  9.210 1.500 9.450 2.460 ;
        RECT  8.930 2.130 9.330 2.530 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.620 2.360 4.380 2.760 ;
        RECT  3.420 2.020 3.860 2.460 ;
        END
    END CP
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.364  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.150 2.740 3.390 ;
        RECT  1.740 3.140 2.180 3.580 ;
        END
    END J
    PIN KZ
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.990 3.060 2.230 ;
        RECT  2.300 1.990 2.740 2.460 ;
        END
    END KZ
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.725  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.250 3.680 18.250 3.920 ;
        RECT  17.420 2.870 18.250 3.920 ;
        RECT  17.700 1.140 17.940 3.920 ;
        RECT  16.220 1.550 17.940 1.790 ;
        RECT  16.220 1.090 16.460 1.790 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.755  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  19.180 1.980 20.900 2.220 ;
        RECT  20.660 1.470 20.900 2.220 ;
        RECT  18.850 3.170 20.560 3.410 ;
        RECT  19.660 3.140 20.100 3.580 ;
        RECT  19.700 1.980 19.940 3.580 ;
        RECT  19.180 1.470 19.420 2.220 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.711  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.910 1.460 13.150 2.480 ;
        RECT  11.100 1.460 13.150 1.700 ;
        RECT  10.750 1.940 11.340 2.180 ;
        RECT  11.100 1.460 11.340 2.180 ;
        RECT  10.420 2.580 11.140 3.020 ;
        RECT  10.750 1.940 10.990 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 21.280 5.600 ;
        RECT  20.720 3.940 21.120 5.600 ;
        RECT  19.410 4.400 19.810 5.600 ;
        RECT  18.110 4.400 18.510 5.600 ;
        RECT  16.740 4.400 17.140 5.600 ;
        RECT  15.200 4.710 15.600 5.600 ;
        RECT  14.270 4.710 14.670 5.600 ;
        RECT  12.830 4.520 13.230 5.600 ;
        RECT  11.440 4.780 11.910 5.600 ;
        RECT  10.070 3.890 10.470 5.600 ;
        RECT  7.840 4.340 8.240 5.600 ;
        RECT  4.240 4.710 4.640 5.600 ;
        RECT  3.380 4.710 3.780 5.600 ;
        RECT  0.880 4.620 1.280 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 21.280 0.740 ;
        RECT  19.840 0.000 20.240 1.610 ;
        RECT  18.360 0.000 18.760 1.350 ;
        RECT  16.880 0.000 17.280 1.210 ;
        RECT  15.130 0.000 15.530 0.890 ;
        RECT  13.920 0.000 14.320 0.890 ;
        RECT  9.310 0.000 9.550 1.260 ;
        RECT  5.050 0.000 5.450 0.890 ;
        RECT  3.940 0.000 4.340 0.890 ;
        RECT  0.890 0.000 1.290 1.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.270 0.470 2.170 ;
        RECT  0.120 1.930 0.900 2.170 ;
        RECT  0.660 1.930 0.900 3.060 ;
        RECT  0.120 1.930 0.360 3.960 ;
        RECT  0.120 3.720 0.690 3.960 ;
        RECT  1.160 1.800 1.400 4.130 ;
        RECT  2.420 3.650 3.350 3.890 ;
        RECT  3.110 3.040 3.350 3.890 ;
        RECT  1.160 3.890 2.660 4.130 ;
        RECT  1.890 0.980 3.540 1.220 ;
        RECT  1.630 1.220 2.130 1.630 ;
        RECT  4.460 1.610 5.040 1.850 ;
        RECT  4.800 1.610 5.040 2.490 ;
        RECT  4.730 2.230 4.970 3.310 ;
        RECT  3.620 3.000 4.300 3.240 ;
        RECT  4.020 3.070 4.970 3.310 ;
        RECT  5.520 1.610 6.220 1.850 ;
        RECT  5.370 2.940 5.760 3.790 ;
        RECT  5.520 1.610 5.760 3.790 ;
        RECT  5.010 3.550 5.760 3.790 ;
        RECT  3.950 1.130 6.920 1.370 ;
        RECT  6.460 1.130 6.920 1.690 ;
        RECT  3.950 1.130 4.190 1.700 ;
        RECT  2.370 1.460 4.190 1.700 ;
        RECT  6.460 1.130 6.700 2.560 ;
        RECT  6.070 2.320 6.700 2.560 ;
        RECT  2.900 4.150 5.670 4.390 ;
        RECT  6.070 2.320 6.310 4.460 ;
        RECT  5.340 4.220 6.310 4.460 ;
        RECT  2.080 4.380 3.140 4.620 ;
        RECT  7.820 1.390 8.400 1.630 ;
        RECT  7.820 1.390 8.060 2.650 ;
        RECT  7.420 2.410 8.060 2.650 ;
        RECT  7.420 2.410 7.660 3.520 ;
        RECT  7.070 3.280 8.830 3.520 ;
        RECT  7.340 1.310 7.580 2.170 ;
        RECT  6.940 1.930 7.580 2.170 ;
        RECT  6.940 1.930 7.180 3.040 ;
        RECT  6.550 2.800 7.180 3.040 ;
        RECT  6.550 3.800 7.570 4.040 ;
        RECT  7.280 3.860 8.720 4.100 ;
        RECT  8.480 3.860 8.720 4.500 ;
        RECT  6.550 2.800 6.790 4.360 ;
        RECT  8.480 4.260 9.370 4.500 ;
        RECT  10.270 1.460 10.860 1.700 ;
        RECT  10.270 1.460 10.510 2.220 ;
        RECT  9.700 1.980 10.510 2.220 ;
        RECT  8.330 2.130 8.570 3.010 ;
        RECT  9.700 1.980 9.940 3.010 ;
        RECT  8.330 2.770 9.940 3.010 ;
        RECT  9.410 3.330 11.070 3.570 ;
        RECT  9.410 2.770 9.650 3.990 ;
        RECT  12.380 2.100 12.620 3.150 ;
        RECT  12.510 2.850 12.750 3.700 ;
        RECT  12.190 3.460 13.510 3.700 ;
        RECT  14.030 2.110 14.270 3.730 ;
        RECT  13.230 3.490 14.270 3.730 ;
        RECT  11.580 1.940 12.140 2.180 ;
        RECT  11.900 1.940 12.140 2.660 ;
        RECT  11.490 2.420 12.140 2.660 ;
        RECT  11.490 2.420 11.730 4.410 ;
        RECT  12.030 3.970 14.750 4.210 ;
        RECT  14.510 2.750 14.750 4.210 ;
        RECT  11.490 4.170 12.290 4.410 ;
        RECT  13.390 1.610 15.230 1.850 ;
        RECT  16.310 2.120 17.330 2.520 ;
        RECT  13.390 1.610 13.630 3.210 ;
        RECT  16.310 2.120 16.550 3.210 ;
        RECT  14.990 2.970 16.550 3.210 ;
        RECT  14.990 1.610 15.230 3.660 ;
    END
END jkbrb4

MACRO jkbrb2
    CLASS CORE ;
    FOREIGN jkbrb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.459  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.540 1.990 16.100 2.390 ;
        RECT  15.820 1.460 16.100 2.390 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.200 2.580 11.700 3.060 ;
        END
    END CP
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.295  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.200 2.360 2.740 3.020 ;
        END
    END J
    PIN KZ
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.840 2.580 4.420 3.020 ;
        END
    END KZ
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.192  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.420 1.460 18.140 1.900 ;
        RECT  17.570 1.460 17.810 3.510 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.192  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.950 1.460 19.440 1.850 ;
        RECT  18.540 3.110 19.190 3.580 ;
        RECT  18.950 1.460 19.190 3.580 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.620 1.460 15.060 1.900 ;
        RECT  14.310 2.710 14.860 3.110 ;
        RECT  14.620 1.460 14.860 3.110 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.160 5.600 ;
        RECT  19.430 4.120 19.670 5.600 ;
        RECT  18.130 4.120 18.370 5.600 ;
        RECT  16.710 4.620 17.110 5.600 ;
        RECT  15.380 4.620 15.780 5.600 ;
        RECT  10.390 4.340 10.630 5.600 ;
        RECT  9.410 4.340 9.650 5.600 ;
        RECT  7.930 4.340 8.170 5.600 ;
        RECT  6.450 4.340 6.690 5.600 ;
        RECT  2.970 4.180 3.210 5.600 ;
        RECT  0.230 3.340 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.160 0.740 ;
        RECT  19.600 0.000 20.000 1.150 ;
        RECT  18.300 0.000 18.700 1.150 ;
        RECT  17.000 0.000 17.400 1.150 ;
        RECT  15.340 0.000 15.580 1.610 ;
        RECT  11.000 0.000 11.240 1.310 ;
        RECT  8.040 0.000 8.280 2.080 ;
        RECT  2.750 0.000 3.150 0.890 ;
        RECT  0.230 0.000 0.470 2.170 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.970 2.730 1.480 3.130 ;
        RECT  0.970 1.770 1.210 3.660 ;
        RECT  2.160 1.130 3.920 1.370 ;
        RECT  2.160 1.130 2.480 1.630 ;
        RECT  1.390 1.010 1.790 1.410 ;
        RECT  4.340 1.240 4.580 1.850 ;
        RECT  2.720 1.610 4.580 1.850 ;
        RECT  1.450 1.010 1.690 2.110 ;
        RECT  2.720 1.610 2.960 2.110 ;
        RECT  1.450 1.870 2.960 2.110 ;
        RECT  1.720 1.870 1.960 4.080 ;
        RECT  1.690 3.680 4.490 3.920 ;
        RECT  1.690 3.680 2.090 4.080 ;
        RECT  4.090 3.680 4.490 4.080 ;
        RECT  5.300 2.090 6.600 2.330 ;
        RECT  5.300 1.480 5.540 3.120 ;
        RECT  4.910 2.880 5.540 3.120 ;
        RECT  4.910 2.880 5.150 4.080 ;
        RECT  5.960 1.560 7.080 1.800 ;
        RECT  6.840 1.560 7.080 2.810 ;
        RECT  6.140 2.570 7.080 2.810 ;
        RECT  6.140 2.570 6.380 4.070 ;
        RECT  5.570 3.830 7.430 4.070 ;
        RECT  7.190 3.830 7.430 4.440 ;
        RECT  10.040 1.460 10.280 2.080 ;
        RECT  9.800 1.840 10.040 3.620 ;
        RECT  11.960 1.460 12.200 2.390 ;
        RECT  10.540 2.050 12.290 2.290 ;
        RECT  11.890 1.990 12.290 2.390 ;
        RECT  10.540 2.050 10.780 3.550 ;
        RECT  10.540 3.310 11.480 3.550 ;
        RECT  12.660 1.460 12.900 2.870 ;
        RECT  11.940 2.630 12.900 2.870 ;
        RECT  6.690 3.120 9.480 3.360 ;
        RECT  9.240 1.480 9.480 4.100 ;
        RECT  9.240 3.860 12.180 4.100 ;
        RECT  11.940 2.630 12.180 4.270 ;
        RECT  11.680 3.860 12.180 4.270 ;
        RECT  8.670 3.120 8.910 4.300 ;
        RECT  8.660 0.980 10.760 1.220 ;
        RECT  11.480 0.980 14.380 1.220 ;
        RECT  4.820 1.000 7.650 1.240 ;
        RECT  10.520 0.980 10.760 1.790 ;
        RECT  11.480 0.980 11.720 1.790 ;
        RECT  10.520 1.550 11.720 1.790 ;
        RECT  7.410 1.000 7.650 2.560 ;
        RECT  4.820 1.000 5.060 2.330 ;
        RECT  3.200 2.090 5.060 2.330 ;
        RECT  14.140 0.980 14.380 2.340 ;
        RECT  13.630 2.100 14.380 2.340 ;
        RECT  8.660 0.980 8.900 2.560 ;
        RECT  7.410 2.320 8.900 2.560 ;
        RECT  3.200 2.090 3.440 3.020 ;
        RECT  13.630 3.390 15.030 3.630 ;
        RECT  13.630 2.100 13.870 3.830 ;
        RECT  13.240 3.590 13.870 3.830 ;
        RECT  13.150 1.460 13.720 1.860 ;
        RECT  13.150 1.460 13.390 3.350 ;
        RECT  12.500 3.110 13.390 3.350 ;
        RECT  15.740 3.110 16.740 3.350 ;
        RECT  12.500 3.110 12.740 4.310 ;
        RECT  15.740 3.110 15.980 4.310 ;
        RECT  12.500 4.070 15.980 4.310 ;
        RECT  16.550 1.430 16.790 2.870 ;
        RECT  16.550 2.140 17.220 2.870 ;
        RECT  15.100 2.630 17.220 2.870 ;
        RECT  15.100 2.630 15.500 3.070 ;
        RECT  16.980 2.140 17.220 3.870 ;
        RECT  16.230 3.630 17.220 3.870 ;
        RECT  16.230 3.630 16.470 4.260 ;
    END
END jkbrb2

MACRO jkbrb1
    CLASS CORE ;
    FOREIGN jkbrb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.020 16.180 2.460 ;
        RECT  15.520 2.220 15.920 2.620 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.210 2.580 11.700 3.060 ;
        END
    END CP
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.295  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.200 2.360 2.740 3.020 ;
        END
    END J
    PIN KZ
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.840 2.580 4.420 3.020 ;
        END
    END KZ
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.108  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.310 3.110 17.860 3.510 ;
        RECT  17.540 1.460 17.860 3.510 ;
        RECT  17.310 1.460 17.860 1.900 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.166  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.540 3.110 19.190 3.580 ;
        RECT  18.950 1.460 19.190 3.580 ;
        RECT  18.790 1.460 19.190 1.850 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.620 2.580 15.060 3.020 ;
        RECT  14.320 2.710 14.720 3.110 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.600 5.600 ;
        RECT  18.130 4.120 18.370 5.600 ;
        RECT  16.790 4.180 17.030 5.600 ;
        RECT  15.460 4.410 15.700 5.600 ;
        RECT  10.390 4.340 10.630 5.600 ;
        RECT  9.410 4.340 9.650 5.600 ;
        RECT  7.930 4.340 8.170 5.600 ;
        RECT  6.450 4.340 6.690 5.600 ;
        RECT  2.970 4.180 3.210 5.600 ;
        RECT  0.230 3.340 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.600 0.740 ;
        RECT  18.130 0.000 18.370 1.330 ;
        RECT  15.350 0.000 15.590 1.830 ;
        RECT  11.010 0.000 11.250 1.310 ;
        RECT  8.050 0.000 8.290 2.080 ;
        RECT  2.760 0.000 3.160 0.890 ;
        RECT  0.230 0.000 0.470 2.170 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.970 2.730 1.480 3.130 ;
        RECT  0.970 1.770 1.210 3.660 ;
        RECT  2.160 1.130 3.930 1.370 ;
        RECT  2.160 1.130 2.480 1.630 ;
        RECT  1.390 1.010 1.790 1.410 ;
        RECT  4.350 1.240 4.590 1.850 ;
        RECT  2.720 1.610 4.590 1.850 ;
        RECT  1.450 1.010 1.690 2.110 ;
        RECT  2.720 1.610 2.960 2.110 ;
        RECT  1.450 1.870 2.960 2.110 ;
        RECT  1.720 1.870 1.960 4.080 ;
        RECT  1.690 3.680 4.490 3.920 ;
        RECT  1.690 3.680 2.090 4.080 ;
        RECT  4.090 3.680 4.490 4.080 ;
        RECT  5.310 2.090 6.610 2.330 ;
        RECT  5.310 1.480 5.550 3.120 ;
        RECT  4.910 2.880 5.550 3.120 ;
        RECT  4.910 2.880 5.150 4.080 ;
        RECT  5.970 1.560 7.090 1.800 ;
        RECT  6.850 1.560 7.090 2.810 ;
        RECT  6.140 2.570 7.090 2.810 ;
        RECT  6.140 2.570 6.380 4.070 ;
        RECT  5.570 3.830 7.430 4.070 ;
        RECT  7.190 3.830 7.430 4.440 ;
        RECT  10.050 1.460 10.290 2.080 ;
        RECT  9.800 1.840 10.290 2.080 ;
        RECT  9.800 1.840 10.040 3.620 ;
        RECT  11.970 1.460 12.210 2.390 ;
        RECT  10.540 2.050 12.290 2.290 ;
        RECT  11.890 1.990 12.290 2.390 ;
        RECT  10.540 2.050 10.780 3.550 ;
        RECT  10.540 3.310 11.480 3.550 ;
        RECT  12.670 1.690 12.910 2.870 ;
        RECT  11.940 2.630 12.910 2.870 ;
        RECT  6.690 3.120 9.490 3.360 ;
        RECT  9.250 1.480 9.490 4.100 ;
        RECT  9.250 3.860 12.180 4.100 ;
        RECT  11.940 2.630 12.180 4.270 ;
        RECT  11.680 3.860 12.180 4.270 ;
        RECT  8.670 3.120 8.910 4.300 ;
        RECT  8.660 0.980 10.770 1.220 ;
        RECT  11.490 0.980 14.390 1.220 ;
        RECT  4.830 1.000 7.650 1.240 ;
        RECT  10.530 0.980 10.770 1.790 ;
        RECT  11.490 0.980 11.730 1.790 ;
        RECT  10.530 1.550 11.730 1.790 ;
        RECT  7.410 1.000 7.650 2.560 ;
        RECT  4.830 1.000 5.070 2.330 ;
        RECT  3.200 2.090 5.070 2.330 ;
        RECT  14.150 0.980 14.390 2.470 ;
        RECT  13.630 2.230 14.390 2.470 ;
        RECT  8.660 0.980 8.900 2.560 ;
        RECT  7.410 2.320 8.900 2.560 ;
        RECT  3.200 2.090 3.440 3.020 ;
        RECT  13.630 3.390 15.030 3.630 ;
        RECT  13.630 2.230 13.870 3.830 ;
        RECT  13.240 3.590 13.870 3.830 ;
        RECT  13.150 1.590 13.730 1.990 ;
        RECT  15.490 2.860 16.560 3.100 ;
        RECT  13.150 1.590 13.390 3.350 ;
        RECT  12.500 3.110 13.390 3.350 ;
        RECT  15.490 2.860 15.730 3.410 ;
        RECT  12.500 3.110 12.740 4.310 ;
        RECT  15.270 3.170 15.510 4.110 ;
        RECT  14.110 3.870 15.510 4.110 ;
        RECT  12.500 4.070 14.350 4.310 ;
        RECT  16.470 1.690 17.040 2.090 ;
        RECT  16.800 2.250 17.300 2.650 ;
        RECT  16.800 1.690 17.040 3.630 ;
        RECT  15.970 3.390 17.040 3.630 ;
    END
END jkbrb1

MACRO invtda
    CLASS CORE ;
    FOREIGN invtda 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.020 1.060 2.460 ;
        RECT  0.600 2.020 0.840 2.880 ;
        END
    END EN
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.660 1.700 9.940 3.020 ;
        RECT  9.540 1.700 9.940 2.100 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.101  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.290 3.460 8.590 4.120 ;
        RECT  8.090 1.210 8.590 4.120 ;
        RECT  4.290 1.210 8.590 1.810 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  8.750 4.350 9.150 5.600 ;
        RECT  7.450 4.350 7.850 5.600 ;
        RECT  6.150 4.350 6.550 5.600 ;
        RECT  4.850 4.350 5.250 5.600 ;
        RECT  3.520 4.710 3.920 5.600 ;
        RECT  0.970 3.900 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  8.750 0.000 9.150 0.980 ;
        RECT  7.450 0.000 7.850 0.980 ;
        RECT  6.150 0.000 6.550 0.980 ;
        RECT  4.850 0.000 5.250 0.980 ;
        RECT  3.550 0.000 3.950 0.980 ;
        RECT  0.890 0.000 1.290 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.140 0.550 1.540 ;
        RECT  0.120 1.140 0.360 4.120 ;
        RECT  1.280 2.740 1.520 3.430 ;
        RECT  0.120 3.190 1.520 3.430 ;
        RECT  0.120 3.190 0.550 4.120 ;
        RECT  1.750 1.770 2.620 2.170 ;
        RECT  3.650 2.830 5.630 3.230 ;
        RECT  1.750 1.770 2.150 4.230 ;
        RECT  1.630 3.670 2.150 4.230 ;
        RECT  3.650 2.830 4.050 4.230 ;
        RECT  1.630 3.830 4.050 4.230 ;
        RECT  2.930 3.830 3.330 4.370 ;
        RECT  1.650 1.130 3.320 1.530 ;
        RECT  2.920 2.050 7.730 2.450 ;
        RECT  2.920 1.130 3.320 3.590 ;
        RECT  2.380 3.190 3.320 3.590 ;
        RECT  8.980 1.220 9.930 1.460 ;
        RECT  8.980 1.220 9.220 3.900 ;
        RECT  8.980 3.660 9.930 3.900 ;
    END
END invtda

MACRO invtd7
    CLASS CORE ;
    FOREIGN invtd7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.140 0.800 2.380 ;
        RECT  0.140 2.140 0.420 3.020 ;
        END
    END EN
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.540 1.700 8.820 3.020 ;
        RECT  8.420 1.700 8.820 2.100 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.825  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.450 3.460 7.450 3.860 ;
        RECT  4.400 1.290 7.400 1.690 ;
        RECT  6.780 1.290 7.220 3.860 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.610 4.350 8.010 5.600 ;
        RECT  6.310 4.350 6.710 5.600 ;
        RECT  5.010 4.350 5.410 5.600 ;
        RECT  3.660 4.440 4.060 5.600 ;
        RECT  0.970 3.900 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.570 0.000 7.970 0.980 ;
        RECT  6.260 0.000 6.660 0.980 ;
        RECT  4.960 0.000 5.360 0.980 ;
        RECT  3.660 0.000 4.060 0.980 ;
        RECT  0.890 0.000 1.290 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.140 0.470 1.900 ;
        RECT  0.230 1.660 1.300 1.900 ;
        RECT  1.060 2.380 2.090 2.620 ;
        RECT  1.060 1.660 1.300 2.870 ;
        RECT  0.810 2.630 1.300 2.870 ;
        RECT  0.810 2.630 1.050 3.620 ;
        RECT  0.230 3.380 1.050 3.620 ;
        RECT  0.230 3.380 0.470 4.120 ;
        RECT  2.220 1.770 2.620 2.170 ;
        RECT  2.380 1.770 2.620 3.100 ;
        RECT  1.710 2.860 2.620 3.100 ;
        RECT  3.970 2.930 5.320 3.170 ;
        RECT  1.710 2.860 1.950 4.060 ;
        RECT  3.970 2.930 4.210 4.060 ;
        RECT  1.710 3.820 4.210 4.060 ;
        RECT  3.000 3.820 3.240 4.620 ;
        RECT  1.650 1.130 3.320 1.370 ;
        RECT  2.920 1.010 3.320 1.600 ;
        RECT  3.070 2.050 6.440 2.290 ;
        RECT  3.070 1.010 3.320 3.580 ;
        RECT  2.380 3.340 3.320 3.580 ;
        RECT  7.860 1.220 8.750 1.460 ;
        RECT  7.860 1.220 8.100 3.900 ;
        RECT  7.860 3.660 8.810 3.900 ;
    END
END invtd7

MACRO invtd4
    CLASS CORE ;
    FOREIGN invtd4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.020 0.800 2.260 ;
        RECT  0.140 2.020 0.420 3.020 ;
        END
    END EN
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.420 1.700 7.700 3.020 ;
        RECT  7.300 1.700 7.700 2.100 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.424  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.590 3.210 6.290 3.450 ;
        RECT  4.390 1.370 6.090 1.610 ;
        RECT  5.100 1.370 5.540 3.450 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  6.450 4.100 6.850 5.600 ;
        RECT  5.030 4.100 5.430 5.600 ;
        RECT  3.660 4.440 4.060 5.600 ;
        RECT  0.970 3.780 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.250 0.000 6.650 0.980 ;
        RECT  4.950 0.000 5.350 0.980 ;
        RECT  3.660 0.000 4.060 0.980 ;
        RECT  0.970 0.000 1.210 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.020 0.470 1.780 ;
        RECT  0.230 1.540 1.300 1.780 ;
        RECT  1.060 2.260 2.090 2.500 ;
        RECT  1.060 1.540 1.300 2.750 ;
        RECT  0.810 2.510 1.300 2.750 ;
        RECT  0.810 2.510 1.050 3.500 ;
        RECT  0.230 3.260 1.050 3.500 ;
        RECT  0.230 3.260 0.470 4.000 ;
        RECT  2.220 1.650 2.620 2.050 ;
        RECT  2.380 1.650 2.620 2.980 ;
        RECT  1.710 2.740 2.620 2.980 ;
        RECT  1.710 2.740 1.950 3.940 ;
        RECT  4.010 2.850 4.250 3.940 ;
        RECT  1.710 3.700 4.250 3.940 ;
        RECT  3.000 3.700 3.240 4.620 ;
        RECT  1.650 1.010 3.310 1.250 ;
        RECT  2.920 1.010 3.310 1.600 ;
        RECT  3.070 1.810 4.250 2.050 ;
        RECT  3.070 1.010 3.310 3.460 ;
        RECT  2.380 3.220 3.310 3.460 ;
        RECT  6.700 1.220 7.570 1.460 ;
        RECT  6.700 1.220 6.940 3.650 ;
        RECT  6.700 3.410 7.650 3.650 ;
    END
END invtd4

MACRO invtd2
    CLASS CORE ;
    FOREIGN invtd2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.640 0.800 3.040 ;
        RECT  0.140 2.640 0.420 3.580 ;
        END
    END EN
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.055  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.580 3.690 2.980 ;
        RECT  2.860 2.580 3.300 3.020 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.310  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.680 2.690 2.080 ;
        RECT  2.380 3.240 2.660 4.140 ;
        RECT  2.280 1.680 2.580 3.640 ;
        RECT  2.250 3.240 2.660 3.640 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  3.370 4.110 3.770 5.600 ;
        RECT  1.050 4.290 1.450 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  3.370 0.000 3.770 1.140 ;
        RECT  0.890 0.000 1.290 1.830 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.640 0.470 2.370 ;
        RECT  0.230 2.130 1.480 2.370 ;
        RECT  1.080 2.130 1.480 3.600 ;
        RECT  0.670 3.360 1.480 3.600 ;
        RECT  0.670 3.360 0.910 4.090 ;
        RECT  0.150 3.850 0.910 4.090 ;
    END
END invtd2

MACRO invtd1
    CLASS CORE ;
    FOREIGN invtd1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.644  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.610 0.800 3.010 ;
        RECT  0.140 2.610 0.420 3.580 ;
        END
    END EN
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.576  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.910 2.020 2.150 3.000 ;
        RECT  1.740 2.020 2.150 2.460 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.568  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.250 4.220 2.660 4.620 ;
        RECT  2.390 0.980 2.660 4.620 ;
        RECT  2.380 3.700 2.660 4.620 ;
        RECT  2.250 0.980 2.660 1.380 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  1.050 4.290 1.450 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  0.890 0.000 1.290 1.830 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.640 0.470 2.370 ;
        RECT  0.230 2.130 1.480 2.370 ;
        RECT  1.080 2.130 1.480 3.570 ;
        RECT  0.740 3.330 1.480 3.570 ;
        RECT  0.740 3.330 0.980 4.060 ;
        RECT  0.150 3.820 0.980 4.060 ;
    END
END invtd1

MACRO invbdk
    CLASS CORE ;
    FOREIGN invbdk 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.998  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.930 1.820 2.330 ;
        RECT  0.480 1.930 1.060 2.460 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 13.775  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.150 2.690 11.640 3.940 ;
        RECT  2.050 1.260 11.640 3.940 ;
        RECT  10.130 1.170 10.530 3.940 ;
        RECT  8.620 1.170 9.020 3.940 ;
        RECT  7.180 1.170 7.580 3.940 ;
        RECT  5.760 1.170 6.160 3.940 ;
        RECT  3.650 1.170 4.050 3.940 ;
        RECT  0.790 1.210 2.590 1.700 ;
        RECT  2.190 1.180 2.590 3.940 ;
        RECT  0.790 1.180 1.190 1.700 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.760 5.600 ;
        RECT  10.330 4.620 10.730 5.600 ;
        RECT  9.000 4.620 9.400 5.600 ;
        RECT  7.670 4.620 8.070 5.600 ;
        RECT  6.340 4.620 6.740 5.600 ;
        RECT  5.010 4.620 5.410 5.600 ;
        RECT  3.400 4.620 3.800 5.600 ;
        RECT  2.070 4.620 2.470 5.600 ;
        RECT  0.740 4.620 1.140 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.760 0.740 ;
        RECT  10.900 0.000 11.300 0.980 ;
        RECT  9.330 0.000 9.730 0.980 ;
        RECT  7.910 0.000 8.310 0.980 ;
        RECT  6.490 0.000 6.890 0.980 ;
        RECT  5.060 0.000 5.460 0.980 ;
        RECT  2.870 0.000 3.270 0.980 ;
        RECT  1.540 0.000 1.940 0.980 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
END invbdk

MACRO invbdf
    CLASS CORE ;
    FOREIGN invbdf 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.470 1.830 1.810 2.230 ;
        RECT  0.470 1.830 1.060 2.460 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 10.956  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.400 1.180 8.840 4.020 ;
        RECT  0.150 2.690 8.840 3.990 ;
        RECT  2.040 1.180 8.840 3.990 ;
        RECT  0.810 1.180 8.840 1.600 ;
        RECT  1.490 2.690 1.890 4.030 ;
        RECT  0.150 2.690 0.550 4.030 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.800 4.620 8.200 5.600 ;
        RECT  6.440 4.620 6.840 5.600 ;
        RECT  5.020 4.230 5.420 5.600 ;
        RECT  3.580 4.230 3.980 5.600 ;
        RECT  2.140 4.620 2.540 5.600 ;
        RECT  0.750 4.620 1.150 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.260 0.000 7.660 0.940 ;
        RECT  5.840 0.000 6.240 0.940 ;
        RECT  4.470 0.000 4.870 0.940 ;
        RECT  2.880 0.000 3.280 0.940 ;
        RECT  1.510 0.000 1.910 0.940 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
END invbdf

MACRO invbda
    CLASS CORE ;
    FOREIGN invbda 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.929  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.480 2.460 1.820 3.020 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.141  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.050 2.580 6.600 3.020 ;
        RECT  5.480 1.220 6.460 4.230 ;
        RECT  5.360 1.060 5.760 3.950 ;
        RECT  0.740 3.310 6.460 3.950 ;
        RECT  2.050 1.220 6.460 3.950 ;
        RECT  3.880 1.060 4.280 3.950 ;
        RECT  2.400 1.060 2.800 3.950 ;
        RECT  0.890 1.220 6.460 1.720 ;
        RECT  0.890 1.040 1.290 1.720 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.410 4.620 5.810 5.600 ;
        RECT  4.080 4.620 4.480 5.600 ;
        RECT  2.780 4.620 3.180 5.600 ;
        RECT  1.480 4.180 1.880 5.600 ;
        RECT  0.150 4.180 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  6.100 0.000 6.500 0.980 ;
        RECT  4.620 0.000 5.020 0.980 ;
        RECT  3.140 0.000 3.540 0.980 ;
        RECT  1.660 0.000 2.060 0.980 ;
        RECT  0.150 0.000 0.550 1.790 ;
        END
    END VSS
END invbda

MACRO invbd7
    CLASS CORE ;
    FOREIGN invbd7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.679  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.110 1.770 4.720 2.170 ;
        RECT  0.410 2.190 2.530 2.590 ;
        RECT  2.110 1.770 2.530 2.590 ;
        RECT  0.620 2.190 1.060 3.020 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.872  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.070 1.220 5.470 2.930 ;
        RECT  0.150 3.540 5.240 3.940 ;
        RECT  4.710 1.020 5.110 1.530 ;
        RECT  4.540 3.140 5.240 3.940 ;
        RECT  4.840 2.690 5.240 3.940 ;
        RECT  1.540 1.220 5.470 1.530 ;
        RECT  3.230 1.020 3.630 1.530 ;
        RECT  1.750 1.020 2.150 1.530 ;
        RECT  0.150 1.660 1.870 1.950 ;
        RECT  1.540 1.220 1.870 1.950 ;
        RECT  0.150 1.020 0.550 1.950 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  3.890 4.620 4.290 5.600 ;
        RECT  2.490 4.620 2.890 5.600 ;
        RECT  0.760 4.180 1.160 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  3.970 0.000 4.370 0.980 ;
        RECT  2.490 0.000 2.890 0.980 ;
        RECT  0.900 0.000 1.300 1.420 ;
        END
    END VSS
END invbd7

MACRO invbd4
    CLASS CORE ;
    FOREIGN invbd4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.318  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.470 2.500 1.060 3.020 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.828  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.920 3.140 3.720 3.540 ;
        RECT  3.200 1.460 3.440 3.540 ;
        RECT  0.360 1.460 3.440 1.890 ;
        RECT  0.720 3.990 2.160 4.230 ;
        RECT  1.920 3.140 2.160 4.230 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  2.660 3.970 2.900 5.600 ;
        RECT  0.150 3.350 1.680 3.610 ;
        RECT  1.280 3.210 1.680 3.610 ;
        RECT  0.150 4.590 0.550 5.600 ;
        RECT  0.150 3.350 0.480 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  2.600 0.000 3.000 1.000 ;
        RECT  0.740 0.000 1.140 1.000 ;
        END
    END VSS
END invbd4

MACRO invbd2
    CLASS CORE ;
    FOREIGN invbd2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.170  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.140 0.870 2.540 ;
        RECT  0.140 2.140 0.500 3.020 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.159  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.740 3.160 2.650 3.450 ;
        RECT  0.150 1.660 2.030 1.900 ;
        RECT  1.630 1.400 2.030 1.900 ;
        RECT  1.180 1.660 1.620 3.450 ;
        RECT  0.150 1.400 0.550 1.900 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  1.760 4.100 2.000 5.600 ;
        RECT  0.230 4.100 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  0.970 0.000 1.210 1.420 ;
        END
    END VSS
END invbd2

MACRO inv0da
    CLASS CORE ;
    FOREIGN inv0da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.590 2.430 1.930 2.830 ;
        RECT  0.590 2.020 1.060 2.830 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.798  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.290 1.700 5.450 3.480 ;
        RECT  3.980 1.700 4.420 3.580 ;
        RECT  1.120 3.060 4.420 3.560 ;
        RECT  1.290 1.700 5.450 2.200 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.560 3.790 4.800 5.600 ;
        RECT  3.250 3.790 3.490 5.600 ;
        RECT  1.940 3.790 2.180 5.600 ;
        RECT  0.550 4.030 0.950 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  5.130 0.000 5.370 1.470 ;
        RECT  3.800 0.000 4.040 1.470 ;
        RECT  2.470 0.000 2.710 1.470 ;
        RECT  1.140 0.000 1.380 1.470 ;
        END
    END VSS
END inv0da

MACRO inv0d7
    CLASS CORE ;
    FOREIGN inv0d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.053  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.500 2.800 2.900 ;
        RECT  0.620 2.500 1.060 3.020 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.972  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.920 3.140 4.530 3.580 ;
        RECT  3.660 1.770 3.940 3.580 ;
        RECT  2.010 1.770 3.940 2.170 ;
        RECT  1.510 3.140 4.530 3.550 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.640 3.990 3.880 5.600 ;
        RECT  2.330 3.990 2.570 5.600 ;
        RECT  0.760 3.450 1.000 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.010 0.000 4.250 1.500 ;
        RECT  2.680 0.000 2.920 1.500 ;
        RECT  1.350 0.000 1.590 1.500 ;
        END
    END VSS
END inv0d7

MACRO inv0d4
    CLASS CORE ;
    FOREIGN inv0d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.922  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.520 0.800 2.920 ;
        RECT  0.140 2.520 0.500 3.580 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.890 3.170 2.620 3.580 ;
        RECT  1.040 3.140 2.620 3.580 ;
        RECT  0.890 1.770 2.620 2.170 ;
        RECT  1.040 1.770 1.320 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.890 3.990 3.130 5.600 ;
        RECT  1.560 3.990 1.800 5.600 ;
        RECT  0.230 3.990 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.890 0.000 3.130 1.500 ;
        RECT  1.560 0.000 1.800 1.500 ;
        RECT  0.230 0.000 0.470 2.100 ;
        END
    END VSS
END inv0d4

MACRO inv0d2
    CLASS CORE ;
    FOREIGN inv0d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.961  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.520 0.800 2.920 ;
        RECT  0.140 2.520 0.500 3.580 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.217  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.890 3.170 1.620 3.580 ;
        RECT  1.040 3.140 1.620 3.580 ;
        RECT  1.040 1.770 1.320 3.580 ;
        RECT  0.890 1.770 1.320 2.170 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.240 5.600 ;
        RECT  1.560 3.990 1.800 5.600 ;
        RECT  0.230 3.990 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.240 0.740 ;
        RECT  1.560 0.000 1.800 1.500 ;
        RECT  0.230 0.000 0.470 2.100 ;
        END
    END VSS
END inv0d2

MACRO inv0d1
    CLASS CORE ;
    FOREIGN inv0d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.520 1.020 2.920 ;
        RECT  0.140 2.520 0.500 3.580 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.110 3.170 1.540 3.570 ;
        RECT  1.260 1.320 1.540 3.570 ;
        RECT  1.110 1.320 1.540 1.720 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 1.680 5.600 ;
        RECT  0.450 3.990 0.690 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 1.680 0.740 ;
        RECT  0.450 0.000 0.690 2.100 ;
        END
    END VSS
END inv0d1

MACRO inv0d0
    CLASS CORE ;
    FOREIGN inv0d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.108  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.790 0.460 3.200 ;
        RECT  0.130 2.510 0.420 3.200 ;
        END
    END I
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.505  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.550 3.430 0.990 3.750 ;
        RECT  0.750 1.740 0.990 3.750 ;
        RECT  0.700 1.740 0.990 2.460 ;
        RECT  0.450 1.740 0.990 2.140 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 1.120 5.600 ;
        RECT  0.440 4.160 0.680 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 1.120 0.740 ;
        RECT  0.430 0.000 0.670 1.340 ;
        END
    END VSS
END inv0d0

MACRO gcnrnna
    CLASS CORE ;
    FOREIGN gcnrnna 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.544  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.930 2.180 2.460 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.420 0.790 2.820 ;
        RECT  0.120 2.420 0.500 3.580 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 7.083  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.120 1.230 8.840 2.960 ;
        RECT  7.720 1.230 8.220 3.450 ;
        RECT  7.590 1.150 7.990 2.960 ;
        RECT  6.100 1.150 6.500 2.960 ;
        RECT  5.220 1.230 5.720 4.320 ;
        RECT  3.180 2.450 5.720 2.980 ;
        RECT  3.140 1.210 5.020 1.590 ;
        RECT  4.620 1.150 5.020 2.980 ;
        RECT  2.710 3.220 3.670 3.720 ;
        RECT  3.180 2.450 3.670 3.720 ;
        RECT  3.140 1.150 3.540 1.590 ;
        END
    END GCLK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  8.480 3.950 8.720 5.600 ;
        RECT  7.000 4.620 7.400 5.600 ;
        RECT  5.700 4.620 6.100 5.600 ;
        RECT  4.660 3.240 4.900 5.600 ;
        RECT  3.360 3.950 3.600 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  8.320 0.000 8.720 0.980 ;
        RECT  6.840 0.000 7.240 0.980 ;
        RECT  5.360 0.000 5.760 0.980 ;
        RECT  3.880 0.000 4.280 0.980 ;
        RECT  2.400 0.000 2.800 0.980 ;
        RECT  0.740 1.090 1.290 1.340 ;
        RECT  0.740 0.000 0.980 1.340 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.040 0.470 2.180 ;
        RECT  0.230 1.940 1.460 2.180 ;
        RECT  1.220 1.630 1.460 4.070 ;
        RECT  0.150 3.830 1.460 4.070 ;
        RECT  1.630 1.030 2.030 1.460 ;
        RECT  1.630 1.220 2.820 1.460 ;
        RECT  2.420 1.820 3.890 2.220 ;
        RECT  2.420 1.220 2.820 2.990 ;
        RECT  2.010 2.690 2.480 3.090 ;
    END
END gcnrnna

MACRO gcnrnn7
    CLASS CORE ;
    FOREIGN gcnrnn7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.546  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.960 2.220 2.460 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.260 0.810 2.660 ;
        RECT  0.120 2.260 0.500 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 4.735  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.200 2.750 6.660 3.150 ;
        RECT  6.220 1.420 6.660 3.150 ;
        RECT  5.990 2.750 6.430 3.490 ;
        RECT  5.990 1.190 6.390 1.660 ;
        RECT  3.030 1.420 6.660 1.660 ;
        RECT  4.510 1.190 4.910 1.660 ;
        RECT  3.030 1.190 3.430 1.660 ;
        END
    END GCLK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.810 4.170 7.050 5.600 ;
        RECT  5.060 4.620 5.460 5.600 ;
        RECT  3.760 4.620 4.160 5.600 ;
        RECT  2.450 4.620 2.850 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.730 0.000 7.130 1.190 ;
        RECT  5.250 0.000 5.650 1.180 ;
        RECT  3.770 0.000 4.170 1.180 ;
        RECT  2.400 0.000 2.800 0.980 ;
        RECT  0.970 0.000 1.210 1.530 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.220 0.470 2.010 ;
        RECT  0.230 1.770 1.460 2.010 ;
        RECT  1.220 1.770 1.460 3.500 ;
        RECT  0.150 3.260 1.460 3.500 ;
        RECT  1.630 1.230 2.700 1.470 ;
        RECT  2.460 1.980 5.850 2.380 ;
        RECT  2.460 1.230 2.700 4.050 ;
        RECT  1.920 3.810 2.700 4.050 ;
    END
END gcnrnn7

MACRO gcnrnn4
    CLASS CORE ;
    FOREIGN gcnrnn4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.549  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.220 2.460 ;
        RECT  1.820 1.880 2.220 2.460 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.460  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.160 0.790 2.560 ;
        RECT  0.120 2.160 0.500 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 3.031  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.470 2.570 6.040 2.970 ;
        RECT  5.660 1.330 6.040 2.970 ;
        RECT  3.220 1.330 6.040 1.570 ;
        RECT  4.700 1.020 4.940 1.570 ;
        RECT  3.220 1.020 3.460 1.570 ;
        END
    END GCLK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.490 4.050 5.730 5.600 ;
        RECT  4.030 4.620 4.430 5.600 ;
        RECT  2.730 4.620 3.130 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.360 0.000 5.760 1.050 ;
        RECT  3.880 0.000 4.280 1.050 ;
        RECT  2.400 0.000 2.800 1.060 ;
        RECT  0.740 1.090 1.290 1.330 ;
        RECT  0.740 0.000 0.980 1.330 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.040 0.470 1.880 ;
        RECT  0.230 1.640 1.480 1.880 ;
        RECT  1.080 1.640 1.480 2.040 ;
        RECT  1.240 1.640 1.480 3.500 ;
        RECT  0.150 3.260 1.480 3.500 ;
        RECT  1.710 1.020 1.950 1.570 ;
        RECT  1.710 1.330 2.700 1.570 ;
        RECT  2.460 1.820 5.420 2.220 ;
        RECT  2.460 1.330 2.700 2.940 ;
        RECT  2.030 2.700 2.700 2.940 ;
    END
END gcnrnn4

MACRO gcnrnn2
    CLASS CORE ;
    FOREIGN gcnrnn2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.553  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.580 1.710 3.020 ;
        RECT  1.470 2.070 1.710 3.020 ;
        RECT  1.160 2.070 1.710 2.310 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.321  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.710 3.020 ;
        RECT  0.470 2.270 0.710 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 1.928  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.360 3.790 4.350 4.030 ;
        RECT  3.980 2.020 4.350 4.030 ;
        RECT  3.450 2.020 4.350 2.260 ;
        RECT  3.450 1.320 3.690 2.260 ;
        RECT  3.270 1.010 3.510 1.560 ;
        END
    END GCLK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.930 4.620 4.330 5.600 ;
        RECT  2.450 4.620 2.860 5.600 ;
        RECT  0.800 3.860 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.930 0.000 4.330 0.980 ;
        RECT  2.420 0.000 2.820 0.890 ;
        RECT  0.740 1.100 1.290 1.340 ;
        RECT  0.740 0.000 0.980 1.340 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.040 0.470 1.830 ;
        RECT  0.230 1.590 2.020 1.830 ;
        RECT  1.860 1.640 2.530 1.880 ;
        RECT  2.290 1.640 2.530 3.500 ;
        RECT  0.150 3.260 2.530 3.500 ;
        RECT  1.650 1.100 2.290 1.340 ;
        RECT  2.160 1.130 3.020 1.370 ;
        RECT  2.780 1.800 3.210 2.200 ;
        RECT  2.780 1.130 3.020 4.030 ;
        RECT  1.420 3.790 3.020 4.030 ;
    END
END gcnrnn2

MACRO gcnrnn1
    CLASS CORE ;
    FOREIGN gcnrnn1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.060 3.020 ;
        RECT  0.620 2.190 0.860 3.020 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.638  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.460 2.250 1.910 ;
        RECT  1.520 1.460 1.760 2.260 ;
        RECT  1.300 1.960 1.560 2.570 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 1.983  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.500 3.740 3.240 3.980 ;
        RECT  2.810 2.100 3.240 3.980 ;
        RECT  2.530 2.100 3.240 2.340 ;
        RECT  2.530 1.400 2.770 2.340 ;
        END
    END GCLK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.810 4.380 3.210 5.600 ;
        RECT  0.740 3.980 1.140 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  0.970 0.000 1.210 1.730 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.140 1.390 0.560 1.820 ;
        RECT  0.140 1.390 0.380 3.660 ;
        RECT  2.010 2.180 2.250 3.500 ;
        RECT  0.140 3.260 2.250 3.500 ;
        RECT  0.140 3.260 0.610 3.660 ;
    END
END gcnrnn1

MACRO gcnfnna
    CLASS CORE ;
    FOREIGN gcnfnna 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.565  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.880 0.550 2.280 ;
        RECT  0.120 1.880 0.500 3.020 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.590  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.860 2.020 1.540 2.460 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 6.914  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.100 1.300 7.240 3.020 ;
        RECT  6.840 1.180 7.240 3.020 ;
        RECT  6.100 1.300 6.600 4.490 ;
        RECT  3.430 1.300 7.240 3.010 ;
        RECT  5.130 0.980 5.370 3.010 ;
        RECT  2.350 1.130 3.890 1.630 ;
        RECT  3.650 0.980 3.890 3.010 ;
        RECT  3.310 2.490 3.820 4.620 ;
        RECT  2.350 2.490 7.240 2.860 ;
        RECT  2.160 3.820 2.600 4.140 ;
        RECT  2.350 2.490 2.600 4.140 ;
        RECT  2.090 0.980 2.590 1.220 ;
        END
    END GCLK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  7.020 3.490 7.420 5.600 ;
        RECT  5.360 3.430 5.760 5.600 ;
        RECT  4.060 3.530 4.460 5.600 ;
        RECT  2.830 3.090 3.070 5.600 ;
        RECT  1.600 4.420 2.000 5.600 ;
        RECT  0.150 3.980 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  5.990 0.000 6.390 0.980 ;
        RECT  4.310 0.000 4.710 0.980 ;
        RECT  2.830 0.000 3.230 0.900 ;
        RECT  1.350 0.000 1.750 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.970 1.120 1.370 ;
        RECT  0.780 0.970 1.120 1.790 ;
        RECT  0.780 1.450 2.110 1.790 ;
        RECT  1.770 1.860 3.200 2.260 ;
        RECT  1.770 1.450 2.110 3.410 ;
        RECT  0.740 2.900 2.110 3.410 ;
    END
END gcnfnna

MACRO gcnfnn7
    CLASS CORE ;
    FOREIGN gcnfnn7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.599  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.100 2.020 1.620 2.460 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.561  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.880 0.630 2.280 ;
        RECT  0.120 1.880 0.500 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 4.641  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.360 6.010 1.600 ;
        RECT  2.830 2.640 5.540 2.880 ;
        RECT  5.100 1.360 5.540 2.880 ;
        RECT  3.580 2.640 3.820 4.320 ;
        RECT  2.200 3.920 3.070 4.160 ;
        RECT  2.830 2.640 3.070 4.160 ;
        END
    END GCLK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.400 4.110 5.800 5.600 ;
        RECT  4.060 3.240 4.460 5.600 ;
        RECT  2.940 4.620 3.340 5.600 ;
        RECT  1.600 4.490 2.000 5.600 ;
        RECT  0.150 3.980 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.530 0.000 4.930 0.980 ;
        RECT  3.220 0.000 3.620 0.980 ;
        RECT  1.880 0.000 2.280 0.890 ;
        RECT  0.150 0.000 0.550 1.010 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.460 1.200 1.700 1.780 ;
        RECT  1.460 1.540 2.100 1.780 ;
        RECT  1.860 1.900 4.420 2.300 ;
        RECT  1.860 1.540 2.100 3.410 ;
        RECT  0.740 3.170 2.100 3.410 ;
    END
END gcnfnn7

MACRO gcnfnn4
    CLASS CORE ;
    FOREIGN gcnfnn4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.553  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.880 0.630 2.280 ;
        RECT  0.120 1.880 0.500 2.460 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.562  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.910 2.580 1.620 3.020 ;
        RECT  0.910 2.030 1.310 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 3.001  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.770 4.420 3.010 ;
        RECT  3.730 2.580 4.420 3.010 ;
        RECT  3.730 1.570 3.970 3.010 ;
        RECT  3.680 1.050 3.920 1.810 ;
        RECT  3.640 2.770 3.880 4.240 ;
        RECT  2.340 1.570 3.970 1.810 ;
        RECT  2.150 3.930 2.580 4.330 ;
        RECT  2.340 2.770 2.580 4.330 ;
        RECT  2.340 0.980 2.580 1.810 ;
        RECT  2.090 0.980 2.580 1.380 ;
        END
    END GCLK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.340 3.840 4.740 5.600 ;
        RECT  2.820 3.250 3.220 5.600 ;
        RECT  1.550 4.620 1.950 5.600 ;
        RECT  0.150 3.980 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.340 0.000 4.740 1.460 ;
        RECT  2.830 0.000 3.230 0.980 ;
        RECT  1.350 0.000 1.750 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.130 1.160 1.370 ;
        RECT  0.920 1.130 1.160 1.780 ;
        RECT  0.920 1.540 1.900 1.780 ;
        RECT  1.660 1.540 1.900 2.320 ;
        RECT  1.860 2.050 3.490 2.450 ;
        RECT  1.860 2.050 2.100 3.600 ;
        RECT  0.740 3.360 2.100 3.600 ;
    END
END gcnfnn4

MACRO gcnfnn2
    CLASS CORE ;
    FOREIGN gcnfnn2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.421  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.790 0.630 2.190 ;
        RECT  0.120 1.790 0.500 3.020 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.433  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.960 2.020 1.620 2.600 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 1.980  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.370 2.220 3.240 2.460 ;
        RECT  2.860 2.020 3.240 2.460 ;
        RECT  2.370 1.480 3.060 1.720 ;
        RECT  2.170 3.910 2.610 4.310 ;
        RECT  2.370 1.480 2.610 4.310 ;
        END
    END GCLK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.890 3.280 3.130 5.600 ;
        RECT  1.620 4.620 2.020 5.600 ;
        RECT  0.150 4.180 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  1.450 0.000 1.850 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.270 2.130 1.510 ;
        RECT  1.890 1.270 2.130 3.080 ;
        RECT  0.800 2.840 2.130 3.080 ;
        RECT  0.800 2.840 1.040 3.830 ;
    END
END gcnfnn2

MACRO gcnfnn1
    CLASS CORE ;
    FOREIGN gcnfnn1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.100 0.800 2.500 ;
        RECT  0.120 2.100 0.500 3.020 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.070 2.520 1.620 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 1.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.390 2.680 1.900 ;
        RECT  2.220 3.730 2.620 4.130 ;
        RECT  2.380 0.990 2.620 4.130 ;
        RECT  2.220 0.990 2.620 1.390 ;
        END
    END GCLK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  1.600 4.560 2.000 5.600 ;
        RECT  0.150 4.180 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  1.450 0.000 1.850 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.270 1.840 1.510 ;
        RECT  1.600 1.270 1.840 2.280 ;
        RECT  1.840 2.040 2.060 2.410 ;
        RECT  1.890 2.180 2.130 3.490 ;
        RECT  1.740 3.250 1.980 3.830 ;
        RECT  0.720 3.590 1.980 3.830 ;
    END
END gcnfnn1

MACRO gclrsna
    CLASS CORE ;
    FOREIGN gclrsna 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.508  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.310 2.020 0.550 2.860 ;
        RECT  0.120 2.020 0.550 2.460 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.350 2.740 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 6.293  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.820 1.210 14.320 4.320 ;
        RECT  10.070 2.880 14.320 3.380 ;
        RECT  11.900 1.210 14.320 3.380 ;
        RECT  12.610 1.210 13.110 4.320 ;
        RECT  10.600 1.210 14.320 1.750 ;
        RECT  11.310 2.880 11.810 4.620 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.540 2.060 6.780 2.830 ;
        RECT  6.220 2.580 6.660 3.020 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.120 5.600 ;
        RECT  14.560 3.260 14.960 5.600 ;
        RECT  13.400 4.620 13.800 5.600 ;
        RECT  12.110 4.620 12.500 5.600 ;
        RECT  10.630 3.680 11.030 5.600 ;
        RECT  9.330 4.320 9.740 5.600 ;
        RECT  8.020 4.340 8.420 5.600 ;
        RECT  6.700 4.250 7.100 5.600 ;
        RECT  4.860 4.350 5.260 5.600 ;
        RECT  2.170 4.110 2.570 5.600 ;
        RECT  0.720 3.740 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.120 0.740 ;
        RECT  14.400 0.000 14.800 0.980 ;
        RECT  12.690 0.000 13.090 0.980 ;
        RECT  11.370 0.000 11.770 0.980 ;
        RECT  10.030 0.000 10.430 0.980 ;
        RECT  6.980 0.000 7.370 1.260 ;
        RECT  4.360 0.000 4.760 0.890 ;
        RECT  1.550 0.000 1.950 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.250 1.750 ;
        RECT  1.010 2.460 1.520 2.860 ;
        RECT  1.010 1.510 1.250 3.370 ;
        RECT  0.150 3.130 1.250 3.370 ;
        RECT  2.800 1.610 3.220 2.010 ;
        RECT  2.980 1.610 3.220 3.860 ;
        RECT  2.770 3.460 3.220 3.860 ;
        RECT  2.180 0.980 4.130 1.220 ;
        RECT  1.590 1.130 2.410 1.370 ;
        RECT  1.590 1.130 1.830 2.220 ;
        RECT  1.760 1.990 2.000 3.520 ;
        RECT  1.490 3.120 2.000 3.520 ;
        RECT  4.100 1.490 4.680 1.730 ;
        RECT  4.100 1.490 4.340 2.410 ;
        RECT  4.010 2.190 4.250 3.390 ;
        RECT  4.010 2.990 4.510 3.390 ;
        RECT  3.620 1.460 3.860 2.000 ;
        RECT  5.260 2.380 5.500 3.070 ;
        RECT  4.940 2.830 5.500 3.070 ;
        RECT  3.460 1.780 3.720 4.410 ;
        RECT  4.940 2.830 5.180 3.870 ;
        RECT  3.460 3.630 5.180 3.870 ;
        RECT  3.460 3.630 3.940 4.410 ;
        RECT  4.920 1.590 6.040 1.910 ;
        RECT  4.820 1.940 5.160 2.120 ;
        RECT  5.720 1.590 6.040 1.990 ;
        RECT  4.920 1.590 5.160 2.120 ;
        RECT  4.580 1.970 5.120 2.180 ;
        RECT  4.580 1.970 5.090 2.210 ;
        RECT  4.580 1.970 4.820 2.590 ;
        RECT  5.740 1.590 5.980 3.290 ;
        RECT  5.710 3.190 5.960 4.060 ;
        RECT  5.420 3.660 5.960 4.060 ;
        RECT  6.170 0.980 6.740 1.220 ;
        RECT  6.500 0.980 6.740 1.740 ;
        RECT  6.500 1.500 7.560 1.740 ;
        RECT  6.950 3.180 7.560 3.420 ;
        RECT  7.320 1.500 7.560 3.420 ;
        RECT  6.200 3.390 7.190 3.640 ;
        RECT  6.200 3.390 6.440 3.960 ;
        RECT  8.250 1.510 8.600 1.910 ;
        RECT  8.250 2.220 9.330 2.460 ;
        RECT  9.090 2.220 9.330 2.780 ;
        RECT  8.250 1.510 8.490 3.900 ;
        RECT  7.460 3.660 8.490 3.900 ;
        RECT  8.830 0.980 9.600 1.380 ;
        RECT  9.200 0.980 9.600 1.850 ;
        RECT  9.570 1.450 9.970 2.380 ;
        RECT  9.570 1.980 11.670 2.380 ;
        RECT  9.570 1.450 9.840 3.460 ;
        RECT  8.840 3.060 9.840 3.460 ;
        RECT  8.840 3.060 9.240 3.850 ;
    END
END gclrsna

MACRO gclrsn7
    CLASS CORE ;
    FOREIGN gclrsn7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.508  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.310 2.020 0.550 2.860 ;
        RECT  0.120 2.020 0.550 2.460 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.350 2.740 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 4.658  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.600 1.270 13.710 1.670 ;
        RECT  10.070 2.980 13.380 3.380 ;
        RECT  12.880 1.270 13.380 3.380 ;
        RECT  12.630 2.980 13.030 4.320 ;
        RECT  11.270 4.380 11.830 4.620 ;
        RECT  11.590 2.980 11.830 4.620 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.540 2.060 6.780 2.830 ;
        RECT  6.220 2.580 6.660 3.020 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 14.000 5.600 ;
        RECT  13.370 4.620 13.770 5.600 ;
        RECT  12.070 4.620 12.470 5.600 ;
        RECT  10.630 3.680 11.030 5.600 ;
        RECT  9.330 4.320 9.740 5.600 ;
        RECT  8.020 4.340 8.420 5.600 ;
        RECT  6.700 4.250 7.100 5.600 ;
        RECT  4.860 4.350 5.260 5.600 ;
        RECT  2.170 4.110 2.570 5.600 ;
        RECT  0.720 3.740 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 14.000 0.740 ;
        RECT  12.710 0.000 13.110 0.980 ;
        RECT  11.340 0.000 11.740 0.980 ;
        RECT  10.030 0.000 10.430 0.980 ;
        RECT  6.980 0.000 7.370 1.260 ;
        RECT  4.360 0.000 4.760 0.890 ;
        RECT  1.550 0.000 1.950 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.250 1.750 ;
        RECT  1.010 2.460 1.520 2.860 ;
        RECT  1.010 1.510 1.250 3.370 ;
        RECT  0.150 3.130 1.250 3.370 ;
        RECT  2.800 1.610 3.220 2.010 ;
        RECT  2.980 1.610 3.220 3.810 ;
        RECT  2.770 3.410 3.220 3.810 ;
        RECT  2.180 0.980 4.130 1.220 ;
        RECT  1.590 1.130 2.410 1.370 ;
        RECT  1.590 1.130 1.830 2.220 ;
        RECT  1.760 1.990 2.000 3.520 ;
        RECT  1.490 3.120 2.000 3.520 ;
        RECT  4.100 1.490 4.680 1.730 ;
        RECT  4.100 1.490 4.340 2.410 ;
        RECT  4.010 2.190 4.250 3.390 ;
        RECT  4.010 2.990 4.510 3.390 ;
        RECT  3.620 1.460 3.860 2.000 ;
        RECT  5.260 2.380 5.500 3.070 ;
        RECT  4.940 2.830 5.500 3.070 ;
        RECT  3.460 1.780 3.720 4.410 ;
        RECT  4.940 2.830 5.180 3.870 ;
        RECT  3.460 3.630 5.180 3.870 ;
        RECT  3.460 3.630 3.940 4.410 ;
        RECT  4.920 1.590 6.040 1.910 ;
        RECT  4.820 1.940 5.160 2.120 ;
        RECT  5.720 1.590 5.980 1.990 ;
        RECT  4.920 1.590 5.160 2.120 ;
        RECT  4.580 1.970 5.120 2.180 ;
        RECT  4.580 1.970 5.090 2.210 ;
        RECT  4.580 1.970 4.820 2.590 ;
        RECT  5.740 1.590 5.980 3.290 ;
        RECT  5.710 3.190 5.960 4.060 ;
        RECT  5.420 3.660 5.960 4.060 ;
        RECT  6.170 0.980 6.740 1.220 ;
        RECT  6.500 0.980 6.740 1.740 ;
        RECT  6.500 1.500 7.560 1.740 ;
        RECT  6.950 3.180 7.560 3.420 ;
        RECT  7.320 1.500 7.560 3.420 ;
        RECT  6.200 3.390 7.190 3.640 ;
        RECT  6.200 3.390 6.440 3.960 ;
        RECT  8.250 1.510 8.600 1.910 ;
        RECT  8.250 2.220 9.330 2.460 ;
        RECT  9.090 2.220 9.330 2.780 ;
        RECT  8.250 1.510 8.490 3.900 ;
        RECT  7.460 3.660 8.490 3.900 ;
        RECT  8.830 0.980 9.440 1.220 ;
        RECT  9.200 0.980 9.440 1.690 ;
        RECT  9.200 1.450 9.810 1.690 ;
        RECT  9.570 1.980 11.200 2.380 ;
        RECT  9.570 1.450 9.810 3.300 ;
        RECT  8.840 3.060 9.810 3.300 ;
        RECT  8.840 3.060 9.080 3.850 ;
    END
END gclrsn7

MACRO gclrsn4
    CLASS CORE ;
    FOREIGN gclrsn4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.508  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.310 2.020 0.550 2.860 ;
        RECT  0.120 2.020 0.550 2.460 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.350 2.740 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 3.047  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.630 1.350 12.430 1.590 ;
        RECT  12.030 1.220 12.430 1.590 ;
        RECT  11.510 2.020 12.260 2.460 ;
        RECT  10.070 3.060 11.910 3.300 ;
        RECT  11.510 1.350 11.910 3.300 ;
        RECT  11.270 4.380 11.830 4.620 ;
        RECT  11.590 1.350 11.830 4.620 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.540 2.060 6.780 2.830 ;
        RECT  6.220 2.580 6.660 3.020 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.880 5.600 ;
        RECT  12.070 4.620 12.470 5.600 ;
        RECT  10.630 3.680 11.030 5.600 ;
        RECT  9.330 4.320 9.740 5.600 ;
        RECT  8.020 4.340 8.420 5.600 ;
        RECT  6.700 4.250 7.100 5.600 ;
        RECT  4.860 4.350 5.260 5.600 ;
        RECT  2.170 4.110 2.570 5.600 ;
        RECT  0.720 3.740 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.880 0.740 ;
        RECT  11.370 0.000 11.770 0.980 ;
        RECT  10.030 0.000 10.430 0.980 ;
        RECT  6.980 0.000 7.370 1.260 ;
        RECT  4.360 0.000 4.760 0.890 ;
        RECT  1.550 0.000 1.950 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.250 1.750 ;
        RECT  1.010 2.460 1.520 2.860 ;
        RECT  1.010 1.510 1.250 3.370 ;
        RECT  0.150 3.130 1.250 3.370 ;
        RECT  2.800 1.610 3.220 2.010 ;
        RECT  2.980 1.610 3.220 3.810 ;
        RECT  2.770 3.410 3.220 3.810 ;
        RECT  2.180 0.980 4.130 1.220 ;
        RECT  1.590 1.130 2.410 1.370 ;
        RECT  1.590 1.130 1.830 2.220 ;
        RECT  1.760 1.990 2.000 3.520 ;
        RECT  1.490 3.120 2.000 3.520 ;
        RECT  4.100 1.490 4.680 1.730 ;
        RECT  4.100 1.490 4.340 2.410 ;
        RECT  4.010 2.190 4.250 3.390 ;
        RECT  4.010 2.990 4.510 3.390 ;
        RECT  3.620 1.460 3.860 2.000 ;
        RECT  5.260 2.380 5.500 3.070 ;
        RECT  4.940 2.830 5.500 3.070 ;
        RECT  3.460 1.780 3.720 4.410 ;
        RECT  4.940 2.830 5.180 3.870 ;
        RECT  3.460 3.630 5.180 3.870 ;
        RECT  3.460 3.630 3.940 4.410 ;
        RECT  4.920 1.590 6.040 1.910 ;
        RECT  4.820 1.940 5.160 2.120 ;
        RECT  5.720 1.590 5.980 1.990 ;
        RECT  4.920 1.590 5.160 2.120 ;
        RECT  4.580 1.970 5.120 2.180 ;
        RECT  4.580 1.970 5.090 2.210 ;
        RECT  4.580 1.970 4.820 2.590 ;
        RECT  5.740 1.590 5.980 3.290 ;
        RECT  5.710 3.190 5.960 4.060 ;
        RECT  5.420 3.660 5.960 4.060 ;
        RECT  6.170 0.980 6.740 1.220 ;
        RECT  6.500 0.980 6.740 1.740 ;
        RECT  6.500 1.500 7.560 1.740 ;
        RECT  6.950 3.180 7.560 3.420 ;
        RECT  7.320 1.500 7.560 3.420 ;
        RECT  6.200 3.390 7.190 3.640 ;
        RECT  6.200 3.390 6.440 3.960 ;
        RECT  8.250 1.510 8.600 1.910 ;
        RECT  8.250 2.220 9.330 2.460 ;
        RECT  9.090 2.220 9.330 2.780 ;
        RECT  8.250 1.510 8.490 3.900 ;
        RECT  7.460 3.660 8.490 3.900 ;
        RECT  8.830 0.980 9.440 1.220 ;
        RECT  9.200 0.980 9.440 1.690 ;
        RECT  9.200 1.450 9.810 1.690 ;
        RECT  9.570 1.980 11.200 2.380 ;
        RECT  9.570 1.450 9.810 3.300 ;
        RECT  8.840 3.060 9.810 3.300 ;
        RECT  8.840 3.060 9.080 3.850 ;
    END
END gclrsn4

MACRO gclrsn2
    CLASS CORE ;
    FOREIGN gclrsn2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.495  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.460 0.760 2.860 ;
        RECT  0.120 2.020 0.500 2.860 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.350 2.740 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 1.682  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.150 3.780 11.080 4.020 ;
        RECT  10.820 1.460 11.080 4.020 ;
        RECT  10.640 1.460 11.080 1.970 ;
        RECT  10.150 3.780 10.390 4.340 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.540 2.060 6.780 2.830 ;
        RECT  6.220 2.580 6.660 3.020 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  10.650 4.620 11.050 5.600 ;
        RECT  9.330 4.320 9.740 5.600 ;
        RECT  7.990 4.400 8.390 5.600 ;
        RECT  6.700 4.340 7.100 5.600 ;
        RECT  4.860 4.350 5.260 5.600 ;
        RECT  2.170 4.110 2.570 5.600 ;
        RECT  0.720 3.740 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  10.080 0.000 10.480 0.980 ;
        RECT  6.980 0.000 7.370 1.260 ;
        RECT  4.360 0.000 4.760 0.890 ;
        RECT  1.550 0.000 1.950 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.250 1.750 ;
        RECT  1.010 2.460 1.520 2.860 ;
        RECT  1.010 1.510 1.250 3.370 ;
        RECT  0.150 3.130 1.250 3.370 ;
        RECT  2.800 1.610 3.220 2.030 ;
        RECT  2.980 1.610 3.220 3.820 ;
        RECT  2.770 3.420 3.220 3.820 ;
        RECT  2.180 0.980 4.130 1.220 ;
        RECT  1.590 1.130 2.410 1.370 ;
        RECT  1.590 1.130 1.830 2.220 ;
        RECT  1.760 1.990 2.000 3.520 ;
        RECT  1.490 3.120 2.000 3.520 ;
        RECT  4.100 1.490 4.680 1.730 ;
        RECT  4.100 1.490 4.340 2.410 ;
        RECT  4.010 2.190 4.250 3.390 ;
        RECT  4.010 2.990 4.510 3.390 ;
        RECT  3.620 1.460 3.860 2.000 ;
        RECT  5.260 2.380 5.500 3.140 ;
        RECT  4.940 2.900 5.500 3.140 ;
        RECT  3.460 1.780 3.720 4.410 ;
        RECT  4.940 2.900 5.180 3.870 ;
        RECT  3.460 3.630 5.180 3.870 ;
        RECT  3.460 3.630 3.940 4.410 ;
        RECT  4.920 1.590 6.040 1.910 ;
        RECT  4.820 1.940 5.160 2.120 ;
        RECT  5.720 1.590 6.040 1.990 ;
        RECT  4.920 1.590 5.160 2.120 ;
        RECT  4.580 1.970 5.120 2.180 ;
        RECT  4.580 1.970 5.090 2.210 ;
        RECT  4.580 1.970 4.900 2.590 ;
        RECT  5.740 1.590 5.980 3.360 ;
        RECT  5.710 3.260 5.960 4.060 ;
        RECT  5.420 3.660 5.960 4.060 ;
        RECT  6.170 0.980 6.740 1.220 ;
        RECT  6.500 0.980 6.740 1.740 ;
        RECT  6.500 1.500 7.560 1.740 ;
        RECT  7.320 1.500 7.560 3.480 ;
        RECT  6.950 3.240 7.560 3.480 ;
        RECT  6.950 3.240 7.190 3.730 ;
        RECT  6.200 3.490 7.190 3.730 ;
        RECT  6.200 3.490 6.440 4.050 ;
        RECT  8.250 1.510 8.600 1.910 ;
        RECT  8.250 2.480 9.540 2.720 ;
        RECT  8.250 1.510 8.490 3.960 ;
        RECT  7.430 3.720 8.490 3.960 ;
        RECT  8.830 0.980 9.440 1.220 ;
        RECT  9.200 0.980 9.440 1.690 ;
        RECT  9.200 1.450 10.310 1.690 ;
        RECT  10.070 1.450 10.310 2.480 ;
        RECT  10.070 2.240 10.580 2.480 ;
        RECT  10.340 2.240 10.580 3.530 ;
        RECT  8.810 3.290 10.580 3.530 ;
        RECT  8.810 3.290 9.050 3.850 ;
    END
END gclrsn2

MACRO gclrsn1
    CLASS CORE ;
    FOREIGN gclrsn1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.478  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.550 3.060 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.326  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.580 3.140 6.100 3.580 ;
        RECT  5.580 2.470 5.820 3.580 ;
        RECT  5.270 2.470 5.820 2.710 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 1.265  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.220 3.130 9.920 3.370 ;
        RECT  9.220 2.580 9.460 3.370 ;
        RECT  9.020 1.260 9.260 3.020 ;
        RECT  8.780 1.260 9.260 1.660 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.419  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.060 1.460 6.660 1.900 ;
        RECT  6.060 1.460 6.300 2.740 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  8.210 4.570 8.610 5.600 ;
        RECT  5.820 4.410 6.060 5.600 ;
        RECT  2.820 4.620 3.220 5.600 ;
        RECT  0.800 4.190 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  9.600 0.000 9.840 1.490 ;
        RECT  7.730 0.000 8.130 0.890 ;
        RECT  5.660 0.000 6.060 0.890 ;
        RECT  2.800 0.000 3.200 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.030 1.750 ;
        RECT  0.790 1.510 1.030 2.260 ;
        RECT  0.790 2.020 1.290 2.260 ;
        RECT  1.050 2.020 1.290 3.060 ;
        RECT  0.790 2.820 1.290 3.060 ;
        RECT  0.790 2.820 1.030 3.540 ;
        RECT  0.150 3.300 1.030 3.540 ;
        RECT  3.570 1.610 4.040 2.010 ;
        RECT  3.800 1.610 4.040 3.420 ;
        RECT  3.530 3.020 4.040 3.420 ;
        RECT  3.430 0.980 4.160 1.220 ;
        RECT  1.510 1.130 3.670 1.370 ;
        RECT  1.510 1.070 1.910 1.470 ;
        RECT  1.530 1.070 1.770 3.840 ;
        RECT  4.420 1.230 4.660 1.750 ;
        RECT  2.490 2.170 2.730 3.340 ;
        RECT  4.310 1.540 4.550 3.900 ;
        RECT  2.710 3.100 2.950 3.900 ;
        RECT  4.280 3.430 4.680 3.900 ;
        RECT  2.710 3.660 4.680 3.900 ;
        RECT  5.160 1.430 5.400 2.230 ;
        RECT  4.790 1.990 5.400 2.230 ;
        RECT  4.790 1.990 5.030 3.190 ;
        RECT  4.790 2.950 5.340 3.190 ;
        RECT  5.100 2.950 5.340 3.580 ;
        RECT  2.010 1.690 3.330 1.930 ;
        RECT  3.090 1.690 3.330 2.460 ;
        RECT  6.540 2.150 7.090 2.550 ;
        RECT  3.200 2.220 3.440 2.780 ;
        RECT  2.010 1.690 2.250 3.820 ;
        RECT  2.230 3.580 2.470 4.380 ;
        RECT  4.960 3.930 6.780 4.170 ;
        RECT  6.540 2.150 6.780 4.170 ;
        RECT  2.230 4.140 5.200 4.380 ;
        RECT  6.900 1.510 7.740 1.750 ;
        RECT  7.500 2.510 8.530 2.750 ;
        RECT  7.020 2.920 7.260 3.500 ;
        RECT  7.500 1.510 7.740 3.500 ;
        RECT  7.020 3.260 7.740 3.500 ;
        RECT  7.470 3.940 10.490 4.180 ;
    END
END gclrsn1

MACRO gclfsna
    CLASS CORE ;
    FOREIGN gclfsna 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.500 2.460 ;
        RECT  0.220 2.020 0.460 2.920 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.348  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.450 2.740 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 7.164  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.140 2.780 15.310 3.260 ;
        RECT  14.900 1.100 15.310 3.260 ;
        RECT  12.420 1.220 15.310 3.260 ;
        RECT  13.420 1.100 13.820 3.260 ;
        RECT  12.360 2.780 12.760 4.580 ;
        RECT  10.410 1.220 15.310 1.620 ;
        RECT  11.940 1.100 12.340 1.620 ;
        RECT  10.410 1.000 10.810 1.620 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 2.010 7.240 2.460 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  15.690 3.700 16.090 5.600 ;
        RECT  14.350 4.270 14.750 5.600 ;
        RECT  13.050 3.490 13.450 5.600 ;
        RECT  11.700 4.610 12.100 5.600 ;
        RECT  10.400 4.270 10.800 5.600 ;
        RECT  7.080 3.180 7.480 5.600 ;
        RECT  4.770 4.360 5.170 5.600 ;
        RECT  2.150 3.260 2.550 5.600 ;
        RECT  0.810 4.410 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  15.640 0.000 16.040 0.980 ;
        RECT  14.160 0.000 14.560 0.980 ;
        RECT  12.680 0.000 13.080 0.980 ;
        RECT  11.200 0.000 11.600 0.980 ;
        RECT  9.340 0.000 9.740 1.380 ;
        RECT  7.810 0.000 8.210 1.290 ;
        RECT  6.270 0.000 6.670 0.890 ;
        RECT  4.980 0.000 5.380 0.890 ;
        RECT  2.230 0.000 2.630 0.900 ;
        RECT  0.740 0.000 1.140 0.900 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.520 1.320 1.760 ;
        RECT  1.080 1.520 1.320 2.910 ;
        RECT  1.080 2.130 1.400 2.910 ;
        RECT  0.970 2.700 1.210 3.710 ;
        RECT  0.150 3.470 1.210 3.710 ;
        RECT  2.980 1.630 3.220 4.030 ;
        RECT  2.800 3.790 3.040 4.360 ;
        RECT  2.960 0.980 3.560 1.220 ;
        RECT  1.600 1.140 3.190 1.380 ;
        RECT  1.600 1.140 1.840 1.980 ;
        RECT  1.640 1.830 1.880 3.780 ;
        RECT  1.450 3.380 1.880 3.780 ;
        RECT  4.290 1.300 4.790 1.700 ;
        RECT  4.290 1.300 4.530 2.230 ;
        RECT  3.940 1.990 4.530 2.230 ;
        RECT  3.940 1.990 4.180 3.490 ;
        RECT  3.940 3.090 4.430 3.490 ;
        RECT  3.460 1.510 4.050 1.750 ;
        RECT  5.400 2.440 5.640 3.440 ;
        RECT  4.760 3.200 5.640 3.440 ;
        RECT  3.460 1.510 3.700 4.000 ;
        RECT  4.760 3.200 5.000 4.000 ;
        RECT  3.460 3.760 5.000 4.000 ;
        RECT  3.540 3.760 3.780 4.620 ;
        RECT  5.340 1.580 6.320 1.820 ;
        RECT  5.340 1.580 5.580 2.180 ;
        RECT  4.770 1.940 5.580 2.180 ;
        RECT  4.770 1.940 5.010 2.710 ;
        RECT  4.420 2.470 5.010 2.710 ;
        RECT  6.080 1.580 6.320 3.920 ;
        RECT  5.350 3.680 6.320 3.920 ;
        RECT  7.120 1.050 7.360 1.770 ;
        RECT  7.120 1.530 7.990 1.770 ;
        RECT  9.310 2.330 9.890 2.570 ;
        RECT  7.750 1.530 7.990 2.940 ;
        RECT  9.310 2.330 9.550 2.940 ;
        RECT  6.560 2.700 9.550 2.940 ;
        RECT  6.560 2.700 6.800 4.620 ;
        RECT  6.050 4.380 6.800 4.620 ;
        RECT  9.130 3.170 10.230 3.410 ;
        RECT  7.820 3.680 9.530 3.920 ;
        RECT  9.130 3.170 9.530 4.000 ;
        RECT  8.550 1.300 8.950 2.090 ;
        RECT  8.550 1.690 10.180 2.090 ;
        RECT  10.120 1.850 12.190 2.250 ;
        RECT  10.480 1.850 10.880 4.040 ;
        RECT  9.760 3.640 10.880 4.040 ;
        RECT  9.760 3.640 10.160 4.630 ;
        RECT  8.390 4.230 10.160 4.630 ;
    END
END gclfsna

MACRO gclfsn7
    CLASS CORE ;
    FOREIGN gclfsn7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.230 2.400 0.630 2.800 ;
        RECT  0.120 2.020 0.500 2.460 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.348  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.350 2.810 2.750 ;
        RECT  2.300 2.350 2.740 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 5.424  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.040 1.240 13.260 1.480 ;
        RECT  12.950 2.360 13.190 3.450 ;
        RECT  9.060 2.360 13.190 2.690 ;
        RECT  11.820 1.240 12.260 2.690 ;
        RECT  11.460 4.380 12.010 4.620 ;
        RECT  11.460 2.360 11.700 4.620 ;
        RECT  10.390 2.360 10.630 4.040 ;
        RECT  9.060 2.360 9.300 3.380 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.580 7.780 3.020 ;
        RECT  7.120 1.860 7.360 2.820 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 13.440 5.600 ;
        RECT  12.350 3.700 12.590 5.600 ;
        RECT  10.950 2.940 11.190 5.600 ;
        RECT  9.750 4.340 10.150 5.600 ;
        RECT  7.070 4.400 7.470 5.600 ;
        RECT  4.770 4.160 5.170 5.600 ;
        RECT  2.120 4.360 2.520 5.600 ;
        RECT  0.720 3.520 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 13.440 0.740 ;
        RECT  12.180 0.000 12.580 0.980 ;
        RECT  10.780 0.000 11.180 0.980 ;
        RECT  9.380 0.000 9.780 0.980 ;
        RECT  7.880 0.000 8.120 1.200 ;
        RECT  6.000 0.000 6.400 0.890 ;
        RECT  5.150 0.000 5.550 0.890 ;
        RECT  2.310 0.000 2.710 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.230 1.750 ;
        RECT  0.990 1.510 1.230 3.280 ;
        RECT  0.230 3.040 1.230 3.280 ;
        RECT  0.230 3.040 0.470 4.620 ;
        RECT  2.900 1.630 3.320 2.030 ;
        RECT  3.080 1.630 3.320 3.730 ;
        RECT  2.690 3.490 3.320 3.730 ;
        RECT  2.990 0.980 3.550 1.220 ;
        RECT  1.590 1.130 3.230 1.370 ;
        RECT  1.590 1.130 1.830 2.680 ;
        RECT  1.500 2.440 1.740 3.360 ;
        RECT  4.200 1.460 4.780 1.700 ;
        RECT  4.200 1.460 4.440 2.410 ;
        RECT  4.110 2.190 4.350 3.390 ;
        RECT  3.720 1.410 3.960 2.000 ;
        RECT  5.380 2.390 5.780 2.840 ;
        RECT  4.710 2.600 5.780 2.840 ;
        RECT  3.560 1.770 3.800 4.410 ;
        RECT  4.710 2.600 4.950 3.870 ;
        RECT  3.560 3.630 4.950 3.870 ;
        RECT  3.560 3.630 3.830 4.410 ;
        RECT  3.430 4.010 3.830 4.410 ;
        RECT  5.020 1.550 6.380 1.790 ;
        RECT  5.020 1.550 5.260 2.180 ;
        RECT  4.680 1.940 5.080 2.360 ;
        RECT  6.140 1.550 6.380 3.320 ;
        RECT  5.340 3.080 6.380 3.320 ;
        RECT  6.640 0.980 7.640 1.220 ;
        RECT  7.400 1.380 7.720 1.620 ;
        RECT  7.400 1.410 7.760 1.620 ;
        RECT  7.400 0.980 7.640 1.620 ;
        RECT  7.480 1.440 8.390 1.650 ;
        RECT  7.520 1.440 8.390 1.680 ;
        RECT  6.640 0.980 6.880 3.810 ;
        RECT  6.040 3.570 6.880 3.810 ;
        RECT  8.570 0.980 9.130 1.220 ;
        RECT  8.890 0.980 9.130 2.120 ;
        RECT  8.580 1.880 11.060 2.120 ;
        RECT  8.890 1.720 11.060 2.120 ;
        RECT  8.350 2.100 8.820 2.340 ;
        RECT  8.350 2.100 8.590 3.920 ;
    END
END gclfsn7

MACRO gclfsn4
    CLASS CORE ;
    FOREIGN gclfsn4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.503  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.320 0.780 2.720 ;
        RECT  0.120 2.320 0.500 3.020 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.348  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.740 3.020 ;
        RECT  2.310 2.260 2.710 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 3.078  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.120 2.020 11.640 2.460 ;
        RECT  11.210 1.170 11.610 1.570 ;
        RECT  9.020 2.410 11.360 2.650 ;
        RECT  11.120 1.250 11.360 2.650 ;
        RECT  9.730 1.250 11.610 1.490 ;
        RECT  10.660 2.410 10.900 4.320 ;
        RECT  9.020 4.180 9.430 4.580 ;
        RECT  9.020 2.410 9.260 4.580 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.300 2.580 7.780 3.020 ;
        RECT  7.300 1.950 7.540 3.020 ;
        RECT  7.000 1.950 7.540 2.350 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.760 5.600 ;
        RECT  11.290 3.050 11.530 5.600 ;
        RECT  9.860 3.480 10.100 5.600 ;
        RECT  9.600 3.480 10.100 3.880 ;
        RECT  7.080 3.370 7.480 5.600 ;
        RECT  4.780 4.160 5.180 5.600 ;
        RECT  2.240 3.280 2.480 5.600 ;
        RECT  0.720 3.920 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.760 0.740 ;
        RECT  10.470 0.000 10.870 0.990 ;
        RECT  8.990 0.000 9.390 1.450 ;
        RECT  6.080 0.000 6.320 1.130 ;
        RECT  1.540 0.000 1.940 0.910 ;
        RECT  0.740 0.000 1.140 1.080 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.700 1.260 1.940 ;
        RECT  1.020 2.140 1.500 2.540 ;
        RECT  1.020 1.700 1.260 3.510 ;
        RECT  0.150 3.270 1.260 3.510 ;
        RECT  2.800 1.700 3.220 2.020 ;
        RECT  2.980 1.700 3.220 4.350 ;
        RECT  2.730 3.950 3.220 4.350 ;
        RECT  2.180 0.980 3.390 1.220 ;
        RECT  2.180 0.980 2.420 1.610 ;
        RECT  1.510 1.370 2.420 1.610 ;
        RECT  1.510 1.370 1.980 1.770 ;
        RECT  1.740 1.370 1.980 4.590 ;
        RECT  1.460 4.190 1.980 4.590 ;
        RECT  4.120 1.640 4.720 1.880 ;
        RECT  4.120 1.640 4.360 3.570 ;
        RECT  3.630 0.980 5.840 1.220 ;
        RECT  3.630 0.980 3.870 4.350 ;
        RECT  3.470 3.950 3.870 4.350 ;
        RECT  5.620 1.630 6.080 2.030 ;
        RECT  4.620 2.130 4.860 2.880 ;
        RECT  5.620 2.460 6.270 2.700 ;
        RECT  5.620 1.630 5.860 2.880 ;
        RECT  4.620 2.640 5.860 2.880 ;
        RECT  5.430 2.640 5.670 3.870 ;
        RECT  6.770 0.990 7.190 1.670 ;
        RECT  6.520 1.430 8.020 1.670 ;
        RECT  7.780 1.430 8.020 2.000 ;
        RECT  6.520 1.430 6.760 4.610 ;
        RECT  6.050 4.370 6.760 4.610 ;
        RECT  8.330 1.690 8.700 1.930 ;
        RECT  8.330 1.050 8.570 1.930 ;
        RECT  8.400 1.930 10.870 2.170 ;
        RECT  8.400 1.690 8.640 4.290 ;
    END
END gclfsn4

MACRO gclfsn2
    CLASS CORE ;
    FOREIGN gclfsn2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.490 0.800 2.890 ;
        RECT  0.120 2.020 0.500 2.890 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.348  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.350 2.740 3.020 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 1.499  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.520 4.030 10.520 4.270 ;
        RECT  10.280 0.980 10.520 4.270 ;
        RECT  10.140 2.580 10.520 3.020 ;
        RECT  10.090 0.980 10.520 1.380 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.442  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 3.140 7.510 3.580 ;
        RECT  7.270 2.590 7.510 3.580 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  10.090 4.620 10.490 5.600 ;
        RECT  8.860 3.770 9.100 5.600 ;
        RECT  7.040 4.620 7.440 5.600 ;
        RECT  4.820 4.170 5.060 5.600 ;
        RECT  2.170 4.370 2.410 5.600 ;
        RECT  0.830 3.690 1.070 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  8.740 0.000 9.140 0.890 ;
        RECT  5.670 0.000 6.070 0.890 ;
        RECT  2.210 0.000 2.610 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.310 1.750 ;
        RECT  1.070 1.510 1.310 2.590 ;
        RECT  1.160 2.350 1.400 3.370 ;
        RECT  0.150 3.130 1.400 3.370 ;
        RECT  2.800 1.630 3.220 2.030 ;
        RECT  2.980 1.630 3.220 3.740 ;
        RECT  2.660 3.500 3.220 3.740 ;
        RECT  4.100 1.460 4.710 1.700 ;
        RECT  4.100 1.460 4.340 2.630 ;
        RECT  4.080 2.390 4.320 3.400 ;
        RECT  3.620 1.630 3.860 2.200 ;
        RECT  5.340 2.390 5.580 2.950 ;
        RECT  4.610 2.710 5.580 2.950 ;
        RECT  3.460 1.960 3.700 4.440 ;
        RECT  4.610 2.710 4.850 3.880 ;
        RECT  3.460 3.640 4.850 3.880 ;
        RECT  3.460 3.640 3.730 4.440 ;
        RECT  4.950 1.610 6.530 1.850 ;
        RECT  4.950 1.610 5.190 2.200 ;
        RECT  4.580 1.960 5.020 2.360 ;
        RECT  6.290 1.610 6.530 2.380 ;
        RECT  5.820 2.140 6.530 2.380 ;
        RECT  5.820 2.140 6.060 3.430 ;
        RECT  5.310 3.190 6.060 3.430 ;
        RECT  2.870 0.980 5.190 1.220 ;
        RECT  6.310 0.980 8.500 1.220 ;
        RECT  1.590 1.130 3.110 1.370 ;
        RECT  4.950 1.130 6.550 1.370 ;
        RECT  1.590 1.130 1.830 2.110 ;
        RECT  1.690 1.870 1.930 4.620 ;
        RECT  1.380 4.380 1.930 4.620 ;
        RECT  6.790 1.520 8.060 1.760 ;
        RECT  7.820 1.520 8.060 2.380 ;
        RECT  7.820 2.140 9.070 2.380 ;
        RECT  6.790 1.520 7.030 2.860 ;
        RECT  6.300 2.620 7.030 2.860 ;
        RECT  6.300 2.620 6.540 4.070 ;
        RECT  6.010 3.670 6.540 4.070 ;
        RECT  8.320 1.520 9.550 1.760 ;
        RECT  9.310 1.520 9.550 2.300 ;
        RECT  9.310 2.060 9.900 2.300 ;
        RECT  7.820 2.780 8.060 3.330 ;
        RECT  9.660 2.060 9.900 3.330 ;
        RECT  7.820 3.090 9.900 3.330 ;
    END
END gclfsn2

MACRO gclfsn1
    CLASS CORE ;
    FOREIGN gclfsn1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.550 0.620 3.020 ;
        END
    END CLK
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.360 2.020 3.860 2.460 ;
        END
    END EN
    PIN GCLK
        DIRECTION OUTPUT ;
        USE CLOCK ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.870 1.240 10.460 1.660 ;
        RECT  10.170 1.240 10.410 4.230 ;
        RECT  8.660 1.680 10.410 1.920 ;
        RECT  9.580 1.460 10.410 1.920 ;
        RECT  8.660 3.030 9.100 3.430 ;
        RECT  8.660 1.680 8.910 3.430 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.484  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.750 3.700 3.310 4.140 ;
        RECT  2.750 2.190 2.990 4.140 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  9.520 4.620 9.920 5.600 ;
        RECT  7.680 4.710 8.080 5.600 ;
        RECT  5.320 4.620 5.720 5.600 ;
        RECT  2.640 4.380 3.040 5.600 ;
        RECT  0.720 4.030 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  8.850 0.000 9.250 1.440 ;
        RECT  6.030 0.000 6.430 0.890 ;
        RECT  2.980 0.000 3.380 1.280 ;
        RECT  0.150 0.000 0.550 1.320 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.720 1.120 1.960 ;
        RECT  0.860 2.540 1.500 2.940 ;
        RECT  0.860 1.720 1.120 3.550 ;
        RECT  0.150 3.310 1.120 3.550 ;
        RECT  1.590 0.980 2.270 1.220 ;
        RECT  1.590 0.980 1.830 2.300 ;
        RECT  1.790 2.060 2.030 3.420 ;
        RECT  1.470 3.180 2.030 3.420 ;
        RECT  4.100 1.460 4.470 1.860 ;
        RECT  4.100 1.460 4.340 2.940 ;
        RECT  3.490 2.700 4.340 2.940 ;
        RECT  3.490 2.700 3.730 3.540 ;
        RECT  5.640 1.660 5.880 2.260 ;
        RECT  5.320 2.020 5.880 2.260 ;
        RECT  5.320 2.020 5.560 3.000 ;
        RECT  5.070 2.760 5.560 3.000 ;
        RECT  5.070 2.760 5.310 3.900 ;
        RECT  4.750 3.660 5.310 3.900 ;
        RECT  4.810 1.460 5.210 1.800 ;
        RECT  4.810 1.460 5.130 1.860 ;
        RECT  4.810 1.460 5.080 2.500 ;
        RECT  4.580 2.260 4.820 3.420 ;
        RECT  4.060 3.180 4.820 3.420 ;
        RECT  6.740 2.530 6.980 3.480 ;
        RECT  5.550 3.240 6.980 3.480 ;
        RECT  4.060 3.180 4.300 4.600 ;
        RECT  4.720 4.140 5.790 4.380 ;
        RECT  5.550 3.240 5.790 4.380 ;
        RECT  4.060 4.360 5.010 4.600 ;
        RECT  6.260 1.690 7.460 1.930 ;
        RECT  6.920 1.660 7.460 2.060 ;
        RECT  6.260 1.690 6.500 2.740 ;
        RECT  5.800 2.500 6.500 2.740 ;
        RECT  7.220 1.660 7.460 3.970 ;
        RECT  6.130 3.720 7.460 3.970 ;
        RECT  6.130 3.720 6.370 4.310 ;
        RECT  3.620 0.980 5.780 1.220 ;
        RECT  6.670 0.980 8.420 1.220 ;
        RECT  5.540 1.130 6.910 1.370 ;
        RECT  3.620 0.980 3.860 1.760 ;
        RECT  2.210 1.520 3.860 1.760 ;
        RECT  2.210 1.520 2.610 1.900 ;
        RECT  2.270 1.520 2.610 1.980 ;
        RECT  8.180 0.980 8.420 2.820 ;
        RECT  2.270 1.520 2.510 4.150 ;
        RECT  2.000 3.760 2.510 4.150 ;
        RECT  9.180 2.190 9.420 2.750 ;
        RECT  7.700 1.460 7.940 3.410 ;
        RECT  7.700 3.090 8.390 3.410 ;
        RECT  8.010 3.090 8.310 3.910 ;
        RECT  9.390 2.510 9.630 3.910 ;
        RECT  8.010 3.670 9.630 3.910 ;
        RECT  8.010 3.090 8.250 4.470 ;
        RECT  6.750 4.230 8.250 4.470 ;
    END
END gclfsn1

MACRO feedth9
    CLASS CORE ;
    FOREIGN feedth9 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        END
    END VSS
END feedth9

MACRO feedth3
    CLASS CORE ;
    FOREIGN feedth3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 1.680 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 1.680 0.740 ;
        END
    END VSS
END feedth3

MACRO feedth
    CLASS CORE ;
    FOREIGN feedth 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 0.560 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 0.560 0.740 ;
        END
    END VSS
END feedth

MACRO dl04d4
    CLASS CORE ;
    FOREIGN dl04d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.433  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.060 3.030 ;
        RECT  0.720 2.200 0.960 3.030 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.051  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.070 1.630 9.790 1.880 ;
        RECT  9.550 1.140 9.790 1.880 ;
        RECT  9.020 2.580 9.460 3.020 ;
        RECT  8.960 3.330 9.360 3.730 ;
        RECT  9.120 1.630 9.360 3.730 ;
        RECT  7.560 3.410 9.360 3.650 ;
        RECT  8.070 1.150 8.310 1.880 ;
        RECT  7.560 3.410 7.800 4.620 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  9.530 4.580 9.930 5.600 ;
        RECT  8.220 3.990 8.630 5.600 ;
        RECT  6.720 4.180 7.120 5.600 ;
        RECT  0.720 4.350 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  8.730 0.000 9.130 1.040 ;
        RECT  7.240 0.000 7.640 1.040 ;
        RECT  0.890 0.000 1.290 1.960 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.130 1.560 0.550 1.960 ;
        RECT  0.130 1.560 0.380 3.760 ;
        RECT  1.680 2.240 1.940 3.600 ;
        RECT  0.130 3.360 1.940 3.600 ;
        RECT  0.130 3.280 0.530 3.760 ;
        RECT  2.270 1.800 3.010 2.060 ;
        RECT  2.770 1.800 3.010 3.460 ;
        RECT  2.500 3.060 3.010 3.460 ;
        RECT  1.550 1.060 3.490 1.300 ;
        RECT  1.550 0.980 1.950 1.380 ;
        RECT  3.250 2.360 4.960 2.600 ;
        RECT  3.250 1.060 3.490 4.500 ;
        RECT  1.420 4.260 3.490 4.500 ;
        RECT  3.750 1.810 5.910 2.050 ;
        RECT  5.670 2.340 6.980 2.580 ;
        RECT  5.670 1.810 5.910 3.360 ;
        RECT  3.730 3.120 5.910 3.360 ;
        RECT  6.620 1.580 7.460 1.820 ;
        RECT  7.220 2.570 8.710 2.810 ;
        RECT  7.220 1.580 7.460 3.060 ;
        RECT  6.310 2.820 7.460 3.060 ;
        RECT  6.310 2.820 6.710 3.280 ;
    END
END dl04d4

MACRO dl04d2
    CLASS CORE ;
    FOREIGN dl04d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.700 1.130 4.140 ;
        RECT  0.730 1.930 1.130 4.140 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.992  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.120 3.050 8.900 3.290 ;
        RECT  8.660 1.300 8.900 3.290 ;
        RECT  8.460 2.580 8.900 3.290 ;
        RECT  8.040 1.300 8.900 1.540 ;
        RECT  8.040 0.990 8.280 1.540 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  8.900 4.080 9.140 5.600 ;
        RECT  7.450 4.620 7.850 5.600 ;
        RECT  3.220 3.840 3.460 5.600 ;
        RECT  0.890 4.620 1.290 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.700 0.000 9.100 0.980 ;
        RECT  7.220 0.000 7.630 0.980 ;
        RECT  5.440 0.000 5.680 1.760 ;
        RECT  0.920 0.000 1.320 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.140 1.730 1.380 ;
        RECT  0.150 1.060 0.550 1.460 ;
        RECT  1.490 1.140 1.730 2.760 ;
        RECT  0.230 1.060 0.470 3.500 ;
        RECT  1.970 1.120 3.190 1.360 ;
        RECT  2.950 1.120 3.190 3.120 ;
        RECT  1.970 1.120 2.210 3.240 ;
        RECT  1.520 3.000 2.210 3.240 ;
        RECT  3.920 2.300 4.160 3.600 ;
        RECT  2.470 3.360 4.160 3.600 ;
        RECT  2.470 1.760 2.710 4.120 ;
        RECT  2.340 3.880 2.580 4.620 ;
        RECT  3.560 1.140 3.800 2.060 ;
        RECT  3.560 1.820 5.200 2.060 ;
        RECT  4.960 1.820 5.200 3.880 ;
        RECT  4.960 3.480 5.600 3.880 ;
        RECT  5.280 3.480 5.520 4.360 ;
        RECT  6.470 2.950 6.710 4.360 ;
        RECT  5.280 4.120 6.710 4.360 ;
        RECT  7.470 1.780 8.410 2.180 ;
        RECT  7.470 1.780 7.790 2.480 ;
        RECT  5.580 2.240 7.790 2.480 ;
        RECT  5.980 2.240 6.220 3.880 ;
    END
END dl04d2

MACRO dl04d1
    CLASS CORE ;
    FOREIGN dl04d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.330 0.720 2.730 ;
        RECT  0.140 2.330 0.500 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.852  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.670 3.210 7.160 3.580 ;
        RECT  6.780 2.580 7.160 3.580 ;
        RECT  6.780 1.460 7.020 3.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.160 4.200 6.400 5.600 ;
        RECT  0.800 4.100 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  5.920 0.000 6.320 0.940 ;
        RECT  1.050 0.000 1.290 1.240 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.400 2.090 ;
        RECT  1.160 1.850 1.400 3.500 ;
        RECT  0.150 3.260 1.400 3.500 ;
        RECT  3.990 1.770 4.230 2.840 ;
        RECT  3.570 2.600 5.570 2.840 ;
        RECT  3.570 2.600 3.810 3.460 ;
        RECT  3.520 0.980 3.930 1.520 ;
        RECT  3.520 1.280 6.470 1.520 ;
        RECT  6.230 1.280 6.470 2.930 ;
        RECT  6.130 2.670 6.370 3.910 ;
        RECT  5.420 3.670 6.370 3.910 ;
        RECT  5.420 3.670 5.660 4.560 ;
        RECT  1.850 4.320 5.660 4.560 ;
    END
END dl04d1

MACRO dl03d4
    CLASS CORE ;
    FOREIGN dl03d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.433  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.880 0.610 2.680 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.780 3.070 7.500 3.580 ;
        RECT  7.260 2.580 7.500 3.580 ;
        RECT  5.290 2.580 7.500 2.820 ;
        RECT  5.070 1.260 6.840 1.500 ;
        RECT  5.290 2.270 5.530 2.820 ;
        RECT  5.070 1.180 5.470 1.580 ;
        RECT  5.070 1.180 5.310 2.510 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.690 4.620 8.090 5.600 ;
        RECT  6.320 4.620 6.720 5.600 ;
        RECT  3.370 3.740 3.770 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.180 0.000 7.580 0.980 ;
        RECT  5.750 0.000 6.160 0.980 ;
        RECT  2.850 0.000 3.250 0.890 ;
        RECT  0.500 0.000 0.900 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.400 1.360 1.640 ;
        RECT  1.120 1.400 1.360 4.130 ;
        RECT  0.150 3.890 1.360 4.130 ;
        RECT  0.150 3.890 0.550 4.290 ;
        RECT  2.240 1.140 2.640 1.540 ;
        RECT  2.240 1.140 2.480 2.850 ;
        RECT  2.910 2.450 3.310 2.850 ;
        RECT  2.080 2.610 3.310 2.850 ;
        RECT  2.080 2.610 2.330 4.080 ;
        RECT  2.080 3.840 2.650 4.080 ;
        RECT  1.620 1.140 1.860 2.020 ;
        RECT  2.890 3.110 4.350 3.350 ;
        RECT  4.110 2.100 4.350 3.770 ;
        RECT  4.110 3.530 4.740 3.770 ;
        RECT  1.600 1.780 1.840 4.620 ;
        RECT  4.500 3.530 4.740 4.490 ;
        RECT  2.890 3.110 3.130 4.620 ;
        RECT  1.600 4.380 3.130 4.620 ;
        RECT  4.300 0.980 4.700 1.860 ;
        RECT  4.590 1.620 4.830 3.290 ;
        RECT  4.590 3.050 5.220 3.290 ;
        RECT  8.120 1.700 8.360 3.550 ;
        RECT  4.980 3.050 5.220 4.130 ;
        RECT  4.980 3.890 5.540 4.130 ;
        RECT  7.880 3.310 8.120 4.380 ;
        RECT  5.300 4.140 8.120 4.380 ;
        RECT  5.300 3.890 5.540 4.610 ;
        RECT  4.980 4.370 5.540 4.610 ;
        RECT  8.190 1.020 8.590 1.420 ;
        RECT  7.820 1.180 8.840 1.420 ;
        RECT  8.190 1.100 8.840 1.420 ;
        RECT  7.350 1.220 8.190 1.460 ;
        RECT  7.350 1.220 7.590 2.030 ;
        RECT  5.600 1.790 7.590 2.030 ;
        RECT  8.600 1.100 8.840 4.190 ;
        RECT  8.390 3.790 8.840 4.190 ;
    END
END dl03d4

MACRO dl03d2
    CLASS CORE ;
    FOREIGN dl03d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.433  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.030 1.060 2.470 ;
        RECT  0.620 2.030 0.860 2.920 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.627  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.530 4.010 7.220 4.250 ;
        RECT  6.980 1.350 7.220 4.250 ;
        RECT  6.780 1.350 7.220 1.900 ;
        RECT  6.240 1.350 7.220 1.590 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  7.100 4.620 7.500 5.600 ;
        RECT  5.790 4.080 6.190 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  5.650 0.000 6.050 0.980 ;
        RECT  0.950 0.000 1.350 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.360 1.780 1.600 ;
        RECT  1.540 1.360 1.780 3.590 ;
        RECT  0.150 3.350 1.780 3.590 ;
        RECT  2.590 1.010 3.180 1.250 ;
        RECT  2.560 1.460 2.830 1.860 ;
        RECT  2.590 1.010 2.830 3.460 ;
        RECT  3.390 1.770 3.630 2.820 ;
        RECT  3.070 2.580 4.380 2.820 ;
        RECT  3.070 2.580 3.310 4.500 ;
        RECT  3.070 4.260 5.100 4.500 ;
        RECT  3.830 0.980 4.480 1.220 ;
        RECT  4.240 0.980 4.480 2.340 ;
        RECT  4.240 2.100 4.860 2.340 ;
        RECT  4.620 2.510 5.400 2.750 ;
        RECT  3.570 3.060 3.810 3.710 ;
        RECT  4.620 2.100 4.860 3.710 ;
        RECT  3.570 3.470 4.860 3.710 ;
        RECT  4.740 1.620 5.900 1.860 ;
        RECT  5.660 1.620 5.900 3.280 ;
        RECT  6.360 2.500 6.600 3.280 ;
        RECT  5.190 3.040 6.600 3.280 ;
    END
END dl03d2

MACRO dl03d1
    CLASS CORE ;
    FOREIGN dl03d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.330 0.720 2.730 ;
        RECT  0.140 2.330 0.500 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.843  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.180 5.480 4.140 ;
        RECT  5.240 1.460 5.480 4.140 ;
        RECT  5.050 1.460 5.480 1.860 ;
        RECT  4.990 3.180 5.480 3.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.490 4.200 4.730 5.600 ;
        RECT  0.800 4.100 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.410 0.000 4.810 0.930 ;
        RECT  1.050 0.000 1.290 1.240 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.400 2.090 ;
        RECT  1.160 1.850 1.400 3.500 ;
        RECT  0.150 3.260 1.400 3.500 ;
        RECT  2.700 1.770 2.940 2.840 ;
        RECT  2.700 2.600 3.890 2.840 ;
        RECT  2.790 2.600 3.030 3.460 ;
        RECT  2.320 0.980 2.730 1.520 ;
        RECT  2.320 1.280 3.990 1.520 ;
        RECT  3.750 1.280 3.990 2.340 ;
        RECT  3.750 2.100 5.000 2.340 ;
        RECT  4.760 2.100 5.000 2.930 ;
        RECT  4.450 2.670 5.000 2.930 ;
        RECT  4.450 2.670 4.690 3.900 ;
        RECT  3.330 3.660 4.690 3.900 ;
        RECT  3.330 3.660 3.620 4.560 ;
        RECT  1.920 4.320 3.620 4.560 ;
    END
END dl03d1

MACRO dl02d4
    CLASS CORE ;
    FOREIGN dl02d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.415  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.460 0.800 2.870 ;
        RECT  0.120 1.810 0.500 2.870 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.831  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.800 1.350 5.560 1.590 ;
        RECT  3.800 4.020 5.420 4.260 ;
        RECT  4.540 1.350 4.980 2.460 ;
        RECT  4.540 1.350 4.780 4.260 ;
        RECT  3.800 3.300 4.040 4.260 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.740 3.050 5.980 5.600 ;
        RECT  5.580 3.050 5.980 3.450 ;
        RECT  4.460 4.620 4.860 5.600 ;
        RECT  3.130 4.710 3.530 5.600 ;
        RECT  0.720 4.370 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.570 0.000 4.970 0.890 ;
        RECT  2.950 0.000 3.340 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.310 1.280 1.550 ;
        RECT  1.040 2.410 1.660 2.810 ;
        RECT  1.040 1.310 1.280 3.370 ;
        RECT  0.150 3.130 1.280 3.370 ;
        RECT  2.530 1.070 2.770 3.980 ;
        RECT  2.530 3.580 3.010 3.980 ;
        RECT  1.790 1.150 2.230 1.550 ;
        RECT  3.250 2.580 3.980 2.820 ;
        RECT  1.990 1.150 2.230 4.470 ;
        RECT  3.250 2.580 3.490 4.470 ;
        RECT  1.480 4.230 3.490 4.470 ;
    END
END dl02d4

MACRO dl02d2
    CLASS CORE ;
    FOREIGN dl02d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.415  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.060 3.020 ;
        RECT  0.720 2.170 0.960 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.552  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.940 2.020 5.480 2.460 ;
        RECT  4.400 2.750 5.180 2.990 ;
        RECT  4.940 1.540 5.180 2.990 ;
        RECT  4.400 2.750 4.640 4.290 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.900 3.230 5.300 5.600 ;
        RECT  3.750 4.620 4.150 5.600 ;
        RECT  0.720 4.520 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.120 0.000 4.520 1.090 ;
        RECT  0.360 0.000 0.760 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.360 1.690 1.640 1.930 ;
        RECT  1.400 1.690 1.640 3.590 ;
        RECT  0.150 3.350 1.640 3.590 ;
        RECT  2.090 1.070 3.070 1.310 ;
        RECT  2.090 1.070 2.330 2.580 ;
        RECT  2.090 2.340 3.170 2.580 ;
        RECT  2.330 2.340 2.570 3.770 ;
        RECT  2.760 1.800 3.650 2.040 ;
        RECT  3.410 2.250 4.690 2.490 ;
        RECT  3.410 1.800 3.650 4.040 ;
        RECT  3.040 3.800 3.650 4.040 ;
        RECT  3.040 3.800 3.280 4.500 ;
        RECT  2.250 4.260 3.280 4.500 ;
    END
END dl02d2

MACRO dl02d1
    CLASS CORE ;
    FOREIGN dl02d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.330 0.720 2.730 ;
        RECT  0.140 2.330 0.500 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.997  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.230 3.180 4.920 3.580 ;
        RECT  4.680 1.460 4.920 3.580 ;
        RECT  4.540 2.480 4.920 3.580 ;
        RECT  4.390 1.460 4.920 1.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.410 4.700 3.810 5.600 ;
        RECT  0.800 4.100 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.620 0.000 4.020 0.940 ;
        RECT  0.980 0.000 1.220 1.240 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.400 2.090 ;
        RECT  1.160 1.850 1.400 3.500 ;
        RECT  0.150 3.260 1.400 3.500 ;
        RECT  2.550 1.770 2.790 2.840 ;
        RECT  2.410 2.600 3.130 2.840 ;
        RECT  2.410 2.600 2.650 3.450 ;
        RECT  2.170 0.980 2.550 1.520 ;
        RECT  2.170 1.280 4.110 1.520 ;
        RECT  3.870 1.280 4.110 2.930 ;
        RECT  3.690 2.670 3.930 4.460 ;
        RECT  1.870 4.220 3.930 4.460 ;
    END
END dl02d1

MACRO dl01d4
    CLASS CORE ;
    FOREIGN dl01d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.800 2.920 ;
        RECT  0.120 2.520 0.420 3.580 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.030 3.020 4.430 3.900 ;
        RECT  2.300 3.020 4.430 3.260 ;
        RECT  2.160 1.230 4.010 1.500 ;
        RECT  3.610 1.100 4.010 1.500 ;
        RECT  2.490 3.020 2.890 3.650 ;
        RECT  2.300 2.580 2.740 3.260 ;
        RECT  2.300 1.230 2.610 3.260 ;
        RECT  2.160 1.100 2.560 1.500 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.610 4.620 5.010 5.600 ;
        RECT  3.230 4.620 3.630 5.600 ;
        RECT  0.720 4.480 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.360 0.000 4.750 0.980 ;
        RECT  2.890 0.000 3.290 0.980 ;
        RECT  0.410 0.000 0.820 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.400 2.090 ;
        RECT  1.160 1.850 1.400 4.120 ;
        RECT  0.150 3.880 1.400 4.120 ;
        RECT  1.440 1.080 1.880 1.480 ;
        RECT  1.640 1.080 1.880 4.580 ;
        RECT  1.640 3.730 2.080 4.580 ;
        RECT  2.620 4.140 6.010 4.380 ;
        RECT  5.610 4.140 6.010 4.480 ;
        RECT  1.640 4.340 2.860 4.580 ;
        RECT  5.000 1.140 6.010 1.380 ;
        RECT  5.000 1.140 5.240 2.140 ;
        RECT  3.140 1.850 5.240 2.140 ;
        RECT  3.140 1.850 4.910 2.250 ;
        RECT  4.670 1.850 4.910 3.840 ;
        RECT  4.670 3.600 5.970 3.840 ;
    END
END dl01d4

MACRO dl01d2
    CLASS CORE ;
    FOREIGN dl01d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.415  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.020 1.060 2.460 ;
        RECT  0.630 2.020 0.870 3.090 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.682  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.890 1.460 4.420 2.010 ;
        RECT  3.990 1.460 4.230 3.560 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.480 4.620 4.880 5.600 ;
        RECT  3.170 4.620 3.570 5.600 ;
        RECT  0.720 4.620 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.080 0.000 3.480 0.910 ;
        RECT  0.950 0.000 1.350 0.910 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.140 1.370 1.640 1.610 ;
        RECT  0.140 1.300 0.550 1.700 ;
        RECT  1.400 1.370 1.640 2.660 ;
        RECT  0.140 1.300 0.380 3.740 ;
        RECT  0.140 3.340 0.550 3.740 ;
        RECT  1.930 2.850 2.920 3.090 ;
        RECT  1.930 2.020 2.170 3.800 ;
        RECT  1.520 3.560 2.170 3.800 ;
        RECT  2.000 1.200 2.930 1.440 ;
        RECT  2.690 1.200 2.930 2.440 ;
        RECT  2.690 2.200 3.740 2.440 ;
        RECT  3.500 2.200 3.740 4.380 ;
        RECT  2.500 4.140 3.740 4.380 ;
    END
END dl01d2

MACRO dl01d1
    CLASS CORE ;
    FOREIGN dl01d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.330 0.720 2.730 ;
        RECT  0.140 2.330 0.500 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.997  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.670 3.130 4.360 3.580 ;
        RECT  4.120 1.460 4.360 3.580 ;
        RECT  3.980 2.480 4.360 3.580 ;
        RECT  3.830 1.460 4.360 1.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  2.850 4.700 3.250 5.600 ;
        RECT  0.800 4.100 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.060 0.000 3.460 0.940 ;
        RECT  0.980 0.000 1.220 1.240 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.400 2.090 ;
        RECT  1.160 1.850 1.400 3.500 ;
        RECT  0.150 3.260 1.400 3.500 ;
        RECT  1.850 1.770 2.100 2.840 ;
        RECT  1.850 2.600 2.570 2.840 ;
        RECT  1.850 1.770 2.090 3.460 ;
        RECT  1.770 0.980 2.170 1.520 ;
        RECT  1.770 1.280 3.470 1.520 ;
        RECT  3.230 1.280 3.470 2.930 ;
        RECT  3.130 2.670 3.370 4.460 ;
        RECT  1.840 4.220 3.370 4.460 ;
    END
END dl01d1

MACRO dfprb4
    CLASS CORE ;
    FOREIGN dfprb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.220 0.780 2.670 ;
        RECT  0.120 2.220 0.500 3.150 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.374  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.170 2.590 2.740 3.130 ;
        RECT  2.170 2.520 2.520 3.130 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.959  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.810 1.960 13.380 2.520 ;
        RECT  12.810 1.160 13.130 2.520 ;
        RECT  11.230 3.120 13.110 3.380 ;
        RECT  12.870 1.160 13.110 3.380 ;
        RECT  11.250 1.420 13.130 1.660 ;
        RECT  12.730 1.160 13.130 1.660 ;
        RECT  11.250 1.160 11.650 1.660 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.000  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.690 1.140 16.050 1.810 ;
        RECT  13.830 3.370 15.940 3.610 ;
        RECT  15.690 1.140 15.930 3.610 ;
        RECT  14.170 1.380 16.050 1.620 ;
        RECT  15.650 1.140 16.050 1.620 ;
        RECT  14.560 3.060 15.120 3.610 ;
        RECT  14.170 1.140 14.570 1.620 ;
        RECT  13.830 3.370 14.230 3.850 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.402  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.300 2.580 5.650 3.110 ;
        RECT  5.100 2.580 5.650 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  15.870 4.360 16.270 5.600 ;
        RECT  14.570 3.990 14.970 5.600 ;
        RECT  13.270 4.180 13.670 5.600 ;
        RECT  11.970 4.170 12.370 5.600 ;
        RECT  10.670 4.130 11.070 5.600 ;
        RECT  8.630 4.710 9.030 5.600 ;
        RECT  5.900 4.430 6.300 5.600 ;
        RECT  4.620 4.610 5.020 5.600 ;
        RECT  1.990 4.100 2.390 5.600 ;
        RECT  0.720 4.090 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  14.910 0.000 15.310 1.020 ;
        RECT  13.430 0.000 13.830 1.030 ;
        RECT  11.990 0.000 12.390 1.010 ;
        RECT  10.510 0.000 10.910 1.360 ;
        RECT  9.620 0.000 10.020 0.890 ;
        RECT  5.000 0.000 5.400 1.750 ;
        RECT  2.010 0.000 2.410 0.890 ;
        RECT  0.440 0.000 0.840 1.070 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.070 1.210 1.670 1.450 ;
        RECT  1.270 1.010 1.670 1.450 ;
        RECT  0.150 1.650 1.260 1.890 ;
        RECT  1.020 1.300 1.260 3.630 ;
        RECT  0.150 3.390 1.260 3.630 ;
        RECT  2.780 1.620 3.250 2.020 ;
        RECT  3.010 1.620 3.250 3.760 ;
        RECT  2.730 3.380 3.250 3.760 ;
        RECT  3.080 0.980 4.150 1.220 ;
        RECT  2.070 1.140 3.320 1.380 ;
        RECT  2.070 1.140 2.310 2.080 ;
        RECT  1.510 1.760 2.310 2.080 ;
        RECT  1.540 1.760 1.910 2.160 ;
        RECT  1.540 1.760 1.780 3.570 ;
        RECT  4.110 1.460 4.660 1.850 ;
        RECT  4.110 1.460 4.350 3.760 ;
        RECT  6.310 2.680 6.550 3.350 ;
        RECT  5.940 3.110 6.550 3.350 ;
        RECT  3.600 4.000 6.180 4.180 ;
        RECT  5.280 3.940 6.180 4.180 ;
        RECT  5.940 3.110 6.180 4.180 ;
        RECT  3.290 4.180 5.520 4.240 ;
        RECT  3.600 1.550 3.840 4.420 ;
        RECT  3.290 4.180 3.840 4.420 ;
        RECT  6.280 1.590 6.520 2.420 ;
        RECT  4.590 2.090 6.520 2.330 ;
        RECT  6.280 2.180 7.030 2.420 ;
        RECT  4.590 2.090 4.830 3.630 ;
        RECT  4.590 3.390 5.700 3.630 ;
        RECT  6.790 2.180 7.030 3.990 ;
        RECT  6.670 3.590 7.030 3.990 ;
        RECT  6.740 1.080 7.990 1.320 ;
        RECT  7.750 1.080 7.990 3.140 ;
        RECT  8.230 1.430 8.470 3.990 ;
        RECT  8.020 3.590 8.470 3.990 ;
        RECT  8.020 3.750 9.800 3.990 ;
        RECT  8.710 1.740 10.760 1.980 ;
        RECT  10.520 1.900 12.460 2.300 ;
        RECT  8.710 1.740 8.950 3.290 ;
        RECT  8.710 3.050 10.330 3.290 ;
        RECT  6.940 1.670 7.510 1.910 ;
        RECT  13.620 1.900 15.350 2.300 ;
        RECT  9.760 2.270 10.160 2.810 ;
        RECT  9.760 2.570 10.810 2.810 ;
        RECT  13.620 1.900 13.860 3.130 ;
        RECT  13.350 2.890 13.860 3.130 ;
        RECT  10.570 2.570 10.810 3.870 ;
        RECT  13.350 2.890 13.590 3.870 ;
        RECT  10.040 3.630 13.590 3.870 ;
        RECT  7.270 1.670 7.510 4.620 ;
        RECT  7.270 4.220 7.700 4.620 ;
        RECT  8.270 4.230 10.280 4.470 ;
        RECT  10.040 3.630 10.280 4.470 ;
        RECT  7.270 4.300 8.450 4.540 ;
        RECT  7.270 4.300 7.800 4.620 ;
    END
END dfprb4

MACRO dfprb2
    CLASS CORE ;
    FOREIGN dfprb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.160 0.790 2.560 ;
        RECT  0.140 2.160 0.500 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.193  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.070 2.100 2.740 2.380 ;
        RECT  2.070 1.820 2.390 2.380 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.318  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.010 3.330 12.820 3.580 ;
        RECT  12.380 3.140 12.820 3.580 ;
        RECT  12.380 1.620 12.620 3.580 ;
        RECT  12.060 1.620 12.620 1.860 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.189  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.440 3.140 14.440 3.650 ;
        RECT  14.050 1.850 14.440 3.650 ;
        RECT  13.440 1.850 14.440 2.090 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.300 2.420 7.010 2.660 ;
        RECT  6.300 1.460 6.690 2.660 ;
        RECT  6.220 1.460 6.690 1.900 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 14.560 5.600 ;
        RECT  14.090 4.280 14.330 5.600 ;
        RECT  12.780 4.290 13.020 5.600 ;
        RECT  11.220 4.710 11.720 5.600 ;
        RECT  9.070 4.650 9.470 5.600 ;
        RECT  6.170 4.710 6.570 5.600 ;
        RECT  4.890 4.700 5.290 5.600 ;
        RECT  2.210 4.620 2.610 5.600 ;
        RECT  0.550 4.200 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 14.560 0.740 ;
        RECT  14.010 0.000 14.410 0.890 ;
        RECT  12.650 0.000 13.050 0.890 ;
        RECT  11.290 0.000 11.690 0.890 ;
        RECT  9.980 0.000 10.220 1.820 ;
        RECT  5.430 0.000 5.670 2.160 ;
        RECT  2.250 0.000 2.650 0.890 ;
        RECT  0.550 0.000 0.790 1.190 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 2.620 2.900 2.860 ;
        RECT  1.590 1.630 1.830 3.600 ;
        RECT  2.860 1.290 3.380 1.610 ;
        RECT  3.140 1.290 3.380 3.820 ;
        RECT  2.800 3.580 3.380 3.820 ;
        RECT  4.420 1.820 4.660 2.730 ;
        RECT  4.360 2.400 4.600 3.900 ;
        RECT  3.620 1.140 4.080 1.580 ;
        RECT  3.620 1.340 5.190 1.580 ;
        RECT  4.950 1.340 5.190 2.660 ;
        RECT  4.950 2.420 6.060 2.660 ;
        RECT  3.620 1.140 3.860 3.900 ;
        RECT  7.050 1.540 7.500 1.940 ;
        RECT  4.910 2.900 5.150 3.570 ;
        RECT  4.910 3.330 7.500 3.570 ;
        RECT  7.260 1.540 7.500 3.800 ;
        RECT  6.940 3.330 7.500 3.800 ;
        RECT  1.030 1.080 2.100 1.320 ;
        RECT  0.150 1.620 1.270 1.860 ;
        RECT  0.150 3.260 1.270 3.500 ;
        RECT  1.030 1.080 1.270 4.260 ;
        RECT  1.030 4.020 2.030 4.260 ;
        RECT  1.770 4.140 4.130 4.380 ;
        RECT  3.730 4.220 7.610 4.460 ;
        RECT  3.730 4.140 4.130 4.600 ;
        RECT  8.600 1.710 8.840 3.130 ;
        RECT  8.530 2.910 8.770 4.230 ;
        RECT  8.530 3.990 10.150 4.230 ;
        RECT  7.780 1.230 9.320 1.470 ;
        RECT  7.780 1.230 8.180 1.960 ;
        RECT  9.080 1.230 9.320 2.530 ;
        RECT  9.080 2.290 10.790 2.530 ;
        RECT  7.780 1.230 8.020 3.800 ;
        RECT  10.640 1.760 11.270 2.000 ;
        RECT  11.030 2.590 12.110 2.830 ;
        RECT  11.030 1.760 11.270 3.010 ;
        RECT  9.650 2.770 11.270 3.010 ;
        RECT  10.530 2.770 10.770 3.760 ;
    END
END dfprb2

MACRO dfprb1
    CLASS CORE ;
    FOREIGN dfprb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.160 0.790 2.560 ;
        RECT  0.140 2.160 0.500 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.193  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.070 2.100 2.740 2.380 ;
        RECT  2.070 1.820 2.390 2.380 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.068  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.580 3.130 12.340 3.580 ;
        RECT  12.100 1.860 12.340 3.580 ;
        RECT  11.590 1.860 12.340 2.100 ;
        RECT  11.590 1.080 11.830 2.100 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.003  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.890 1.560 13.320 3.450 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.300 2.420 7.010 2.660 ;
        RECT  6.300 1.460 6.690 2.660 ;
        RECT  6.220 1.460 6.690 1.900 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 13.440 5.600 ;
        RECT  12.400 4.030 12.640 5.600 ;
        RECT  11.030 4.580 11.430 5.600 ;
        RECT  9.070 4.650 9.470 5.600 ;
        RECT  6.170 4.710 6.570 5.600 ;
        RECT  4.890 4.700 5.290 5.600 ;
        RECT  2.210 4.620 2.610 5.600 ;
        RECT  0.550 4.200 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 13.440 0.740 ;
        RECT  12.290 0.000 12.690 0.890 ;
        RECT  9.980 0.000 10.220 1.820 ;
        RECT  5.430 0.000 5.670 2.160 ;
        RECT  2.250 0.000 2.650 0.890 ;
        RECT  0.550 0.000 0.790 1.190 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 2.620 2.900 2.860 ;
        RECT  1.590 1.630 1.830 3.600 ;
        RECT  2.860 1.290 3.380 1.610 ;
        RECT  3.140 1.290 3.380 3.820 ;
        RECT  2.800 3.580 3.380 3.820 ;
        RECT  4.420 1.820 4.660 2.730 ;
        RECT  4.360 2.400 4.600 3.900 ;
        RECT  3.620 1.140 4.080 1.580 ;
        RECT  3.620 1.340 5.190 1.580 ;
        RECT  4.950 1.340 5.190 2.660 ;
        RECT  4.950 2.420 6.060 2.660 ;
        RECT  3.620 1.140 3.860 3.900 ;
        RECT  7.050 1.540 7.500 1.940 ;
        RECT  4.910 2.900 5.150 3.570 ;
        RECT  4.910 3.330 7.500 3.570 ;
        RECT  7.260 1.540 7.500 3.800 ;
        RECT  6.950 3.330 7.500 3.800 ;
        RECT  1.030 1.080 2.100 1.320 ;
        RECT  0.150 1.620 1.270 1.860 ;
        RECT  0.150 3.260 1.270 3.500 ;
        RECT  1.030 1.080 1.270 4.260 ;
        RECT  1.030 4.020 2.030 4.260 ;
        RECT  1.770 4.140 4.130 4.380 ;
        RECT  3.730 4.220 7.610 4.460 ;
        RECT  3.730 4.140 4.130 4.600 ;
        RECT  8.600 1.710 8.840 3.130 ;
        RECT  8.530 2.910 8.770 4.230 ;
        RECT  8.530 3.990 10.150 4.230 ;
        RECT  7.780 1.230 9.320 1.470 ;
        RECT  7.780 1.230 8.180 1.960 ;
        RECT  9.080 1.230 9.320 2.530 ;
        RECT  9.080 2.290 10.790 2.530 ;
        RECT  7.780 1.230 8.020 3.800 ;
        RECT  10.640 1.760 11.270 2.000 ;
        RECT  11.030 2.590 11.860 2.830 ;
        RECT  11.030 1.760 11.270 3.010 ;
        RECT  9.650 2.770 11.270 3.010 ;
        RECT  10.360 2.770 10.600 3.620 ;
    END
END dfprb1

MACRO dfpfb4
    CLASS CORE ;
    FOREIGN dfpfb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.630 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.180 2.310 2.740 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.890  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.540 3.670 13.380 3.910 ;
        RECT  12.940 1.740 13.380 3.910 ;
        RECT  12.880 1.010 13.280 2.080 ;
        RECT  12.840 3.470 13.380 3.910 ;
        RECT  11.680 1.840 13.380 2.080 ;
        RECT  11.680 1.090 11.920 2.080 ;
        RECT  11.340 1.090 11.920 1.330 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.961  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.850 1.730 16.570 1.970 ;
        RECT  16.330 1.090 16.570 1.970 ;
        RECT  15.440 3.070 15.840 3.470 ;
        RECT  15.180 1.730 15.620 3.390 ;
        RECT  14.140 3.150 15.840 3.390 ;
        RECT  14.850 1.090 15.090 1.970 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.360 2.450 6.100 3.030 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  16.180 4.400 16.580 5.600 ;
        RECT  14.880 4.400 15.280 5.600 ;
        RECT  13.580 4.400 13.980 5.600 ;
        RECT  12.280 4.400 12.680 5.600 ;
        RECT  10.980 4.360 11.380 5.600 ;
        RECT  9.020 4.710 9.430 5.600 ;
        RECT  6.250 4.340 6.650 5.600 ;
        RECT  4.710 4.340 5.110 5.600 ;
        RECT  1.970 4.710 2.380 5.600 ;
        RECT  0.800 4.150 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  15.510 0.000 15.910 0.980 ;
        RECT  13.950 0.000 14.350 1.070 ;
        RECT  12.110 0.000 12.510 0.940 ;
        RECT  10.550 0.000 10.950 0.890 ;
        RECT  9.320 0.000 9.730 0.890 ;
        RECT  4.860 0.000 5.270 0.890 ;
        RECT  2.430 0.000 2.840 0.890 ;
        RECT  0.240 0.000 0.650 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.350 0.980 1.590 1.530 ;
        RECT  0.960 1.290 1.590 1.530 ;
        RECT  0.150 1.750 1.200 1.990 ;
        RECT  0.960 1.290 1.200 3.500 ;
        RECT  0.150 3.260 1.200 3.500 ;
        RECT  2.800 1.670 3.220 2.070 ;
        RECT  2.980 1.670 3.220 4.210 ;
        RECT  2.750 3.810 3.220 4.210 ;
        RECT  3.120 0.980 3.520 1.380 ;
        RECT  1.830 1.140 3.520 1.380 ;
        RECT  1.830 1.140 2.070 2.080 ;
        RECT  1.510 1.770 2.070 2.080 ;
        RECT  1.590 1.770 1.830 3.050 ;
        RECT  1.540 2.740 1.780 3.710 ;
        RECT  4.200 1.630 4.680 2.030 ;
        RECT  4.200 1.630 4.440 3.550 ;
        RECT  3.460 1.620 3.940 2.020 ;
        RECT  6.340 2.540 6.740 2.940 ;
        RECT  6.340 2.540 6.580 3.620 ;
        RECT  4.780 3.380 6.580 3.620 ;
        RECT  3.460 1.620 3.700 4.100 ;
        RECT  4.780 3.380 5.030 4.100 ;
        RECT  3.460 3.860 5.030 4.100 ;
        RECT  3.860 0.980 4.260 1.380 ;
        RECT  5.530 0.980 7.090 1.220 ;
        RECT  3.860 1.140 5.790 1.380 ;
        RECT  6.310 1.500 6.860 1.910 ;
        RECT  4.920 1.670 6.860 1.910 ;
        RECT  6.620 1.500 6.860 2.250 ;
        RECT  6.620 2.010 7.250 2.250 ;
        RECT  4.920 1.670 5.160 2.310 ;
        RECT  4.880 2.170 5.120 2.750 ;
        RECT  4.680 2.350 5.120 2.750 ;
        RECT  7.010 2.010 7.250 4.100 ;
        RECT  5.480 3.860 7.250 4.100 ;
        RECT  8.090 1.460 8.330 2.050 ;
        RECT  8.230 1.810 8.470 3.520 ;
        RECT  8.230 3.280 10.110 3.520 ;
        RECT  7.610 0.980 9.020 1.220 ;
        RECT  8.780 1.130 10.580 1.370 ;
        RECT  7.100 1.530 7.850 1.770 ;
        RECT  10.340 1.130 10.580 2.560 ;
        RECT  10.340 2.160 10.740 2.560 ;
        RECT  7.610 0.980 7.850 2.590 ;
        RECT  7.750 2.310 7.990 3.790 ;
        RECT  8.720 2.540 10.090 2.780 ;
        RECT  9.850 1.630 10.090 3.040 ;
        RECT  8.720 2.540 9.120 2.940 ;
        RECT  11.170 1.660 11.410 3.040 ;
        RECT  9.850 2.800 11.410 3.040 ;
        RECT  10.440 2.800 10.680 4.410 ;
        RECT  10.240 4.010 10.680 4.410 ;
    END
END dfpfb4

MACRO dfpfb2
    CLASS CORE ;
    FOREIGN dfpfb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.160 0.790 2.560 ;
        RECT  0.140 2.160 0.500 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.193  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.460 2.700 2.220 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.318  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.010 3.330 12.820 3.580 ;
        RECT  12.380 3.140 12.820 3.580 ;
        RECT  12.380 1.620 12.620 3.580 ;
        RECT  12.060 1.620 12.620 1.860 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.189  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.440 3.140 14.440 3.650 ;
        RECT  14.050 1.850 14.440 3.650 ;
        RECT  13.440 1.850 14.440 2.090 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.300 2.420 7.010 2.660 ;
        RECT  6.300 1.460 6.690 2.660 ;
        RECT  6.220 1.460 6.690 1.900 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 14.560 5.600 ;
        RECT  14.090 4.280 14.330 5.600 ;
        RECT  12.780 4.290 13.020 5.600 ;
        RECT  11.220 4.710 11.720 5.600 ;
        RECT  9.070 4.650 9.470 5.600 ;
        RECT  6.170 4.710 6.570 5.600 ;
        RECT  4.890 4.700 5.290 5.600 ;
        RECT  2.290 4.380 2.530 5.600 ;
        RECT  0.550 4.200 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 14.560 0.740 ;
        RECT  14.010 0.000 14.410 0.890 ;
        RECT  12.650 0.000 13.050 0.890 ;
        RECT  11.290 0.000 11.690 0.890 ;
        RECT  9.980 0.000 10.220 1.820 ;
        RECT  5.430 0.000 5.670 2.160 ;
        RECT  2.250 0.000 2.650 0.890 ;
        RECT  0.820 0.000 1.060 1.190 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.620 1.270 1.860 ;
        RECT  0.150 3.260 1.270 3.500 ;
        RECT  1.030 1.620 1.270 4.260 ;
        RECT  1.030 4.020 1.670 4.260 ;
        RECT  2.940 1.290 3.180 3.130 ;
        RECT  2.880 2.880 3.120 3.660 ;
        RECT  4.420 1.820 4.660 2.730 ;
        RECT  4.360 2.400 4.600 3.830 ;
        RECT  3.620 1.140 4.080 1.580 ;
        RECT  3.620 1.340 5.190 1.580 ;
        RECT  4.950 1.340 5.190 2.660 ;
        RECT  4.950 2.420 6.060 2.660 ;
        RECT  3.620 1.140 3.860 3.660 ;
        RECT  7.040 1.540 7.490 1.940 ;
        RECT  4.910 2.900 5.150 3.570 ;
        RECT  4.910 3.330 7.490 3.570 ;
        RECT  7.250 1.540 7.490 3.800 ;
        RECT  6.940 3.330 7.490 3.800 ;
        RECT  1.510 1.080 2.100 1.320 ;
        RECT  1.510 1.080 1.770 3.780 ;
        RECT  1.510 1.630 1.910 3.780 ;
        RECT  1.910 3.540 2.150 4.140 ;
        RECT  1.910 3.900 4.130 4.140 ;
        RECT  3.730 3.900 4.130 4.460 ;
        RECT  3.730 4.220 7.610 4.460 ;
        RECT  8.600 1.710 8.840 3.130 ;
        RECT  8.530 2.910 8.770 4.230 ;
        RECT  8.530 3.990 10.150 4.230 ;
        RECT  7.780 1.230 9.320 1.470 ;
        RECT  7.780 1.230 8.180 1.960 ;
        RECT  9.080 1.230 9.320 2.530 ;
        RECT  9.080 2.290 10.790 2.530 ;
        RECT  7.780 1.230 8.020 3.800 ;
        RECT  10.640 1.760 11.270 2.000 ;
        RECT  11.030 2.590 12.110 2.830 ;
        RECT  11.030 1.760 11.270 3.010 ;
        RECT  9.650 2.770 11.270 3.010 ;
        RECT  10.530 2.770 10.770 3.760 ;
    END
END dfpfb2

MACRO dfpfb1
    CLASS CORE ;
    FOREIGN dfpfb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.160 0.790 2.560 ;
        RECT  0.140 2.160 0.500 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.193  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.460 2.700 2.220 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.068  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.580 3.130 12.340 3.580 ;
        RECT  12.100 1.860 12.340 3.580 ;
        RECT  11.590 1.860 12.340 2.100 ;
        RECT  11.590 1.080 11.830 2.100 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.003  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.890 1.560 13.320 3.450 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.300 2.420 7.010 2.660 ;
        RECT  6.300 1.460 6.690 2.660 ;
        RECT  6.220 1.460 6.690 1.900 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 13.440 5.600 ;
        RECT  12.400 4.030 12.640 5.600 ;
        RECT  11.030 4.580 11.430 5.600 ;
        RECT  9.070 4.650 9.470 5.600 ;
        RECT  6.170 4.710 6.570 5.600 ;
        RECT  4.890 4.700 5.290 5.600 ;
        RECT  2.290 4.380 2.530 5.600 ;
        RECT  0.550 4.200 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 13.440 0.740 ;
        RECT  12.290 0.000 12.690 0.890 ;
        RECT  9.980 0.000 10.220 1.820 ;
        RECT  5.430 0.000 5.670 2.160 ;
        RECT  2.250 0.000 2.650 0.890 ;
        RECT  0.820 0.000 1.060 1.190 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.620 1.270 1.860 ;
        RECT  0.150 3.260 1.270 3.500 ;
        RECT  1.030 1.620 1.270 4.260 ;
        RECT  1.030 4.020 1.670 4.260 ;
        RECT  2.940 1.290 3.180 3.130 ;
        RECT  2.880 2.880 3.120 3.660 ;
        RECT  4.420 1.820 4.660 2.730 ;
        RECT  4.360 2.400 4.600 3.830 ;
        RECT  3.620 1.140 4.080 1.580 ;
        RECT  3.620 1.340 5.190 1.580 ;
        RECT  4.950 1.340 5.190 2.660 ;
        RECT  4.950 2.420 6.060 2.660 ;
        RECT  3.620 1.140 3.860 3.660 ;
        RECT  7.040 1.540 7.490 1.940 ;
        RECT  4.910 2.900 5.150 3.570 ;
        RECT  4.910 3.330 7.490 3.570 ;
        RECT  7.250 1.540 7.490 3.800 ;
        RECT  6.940 3.330 7.490 3.800 ;
        RECT  1.510 1.080 2.100 1.320 ;
        RECT  1.510 1.080 1.770 3.780 ;
        RECT  1.510 1.630 1.910 3.780 ;
        RECT  1.910 3.540 2.150 4.140 ;
        RECT  1.910 3.900 4.130 4.140 ;
        RECT  3.730 3.900 4.130 4.460 ;
        RECT  3.730 4.220 7.610 4.460 ;
        RECT  8.600 1.710 8.840 3.130 ;
        RECT  8.530 2.910 8.770 4.230 ;
        RECT  8.530 3.990 10.150 4.230 ;
        RECT  7.780 1.230 9.320 1.470 ;
        RECT  7.780 1.230 8.180 1.960 ;
        RECT  9.080 1.230 9.320 2.530 ;
        RECT  9.080 2.290 10.790 2.530 ;
        RECT  7.780 1.230 8.020 3.800 ;
        RECT  10.640 1.760 11.270 2.000 ;
        RECT  11.030 2.590 11.860 2.830 ;
        RECT  11.030 1.760 11.270 3.010 ;
        RECT  9.650 2.770 11.270 3.010 ;
        RECT  10.360 2.770 10.600 3.620 ;
    END
END dfpfb1

MACRO dfnrq4
    CLASS CORE ;
    FOREIGN dfnrq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.810 2.700 ;
        RECT  0.120 2.300 0.500 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.380  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.160 2.510 2.740 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.062  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.600 3.190 12.200 3.430 ;
        RECT  11.820 1.680 12.200 3.430 ;
        RECT  9.480 1.680 12.200 1.920 ;
        RECT  9.600 2.980 10.000 3.430 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.320 5.600 ;
        RECT  11.480 4.620 11.880 5.600 ;
        RECT  10.160 3.680 10.560 5.600 ;
        RECT  8.860 4.450 9.260 5.600 ;
        RECT  7.590 4.440 7.990 5.600 ;
        RECT  5.180 4.380 5.420 5.600 ;
        RECT  4.770 4.380 5.420 4.620 ;
        RECT  2.140 4.710 2.540 5.600 ;
        RECT  0.720 3.870 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.320 0.740 ;
        RECT  11.530 1.120 12.100 1.360 ;
        RECT  11.530 0.000 11.770 1.360 ;
        RECT  10.220 1.170 10.800 1.420 ;
        RECT  10.560 0.000 10.800 1.420 ;
        RECT  8.040 0.000 8.440 1.520 ;
        RECT  5.050 0.000 5.450 1.680 ;
        RECT  2.140 0.000 2.540 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.490 0.470 2.060 ;
        RECT  0.230 1.820 1.290 2.060 ;
        RECT  1.050 1.820 1.290 2.370 ;
        RECT  1.170 2.130 1.410 3.500 ;
        RECT  0.160 3.260 1.410 3.500 ;
        RECT  2.800 1.690 3.310 2.090 ;
        RECT  3.070 1.690 3.310 3.690 ;
        RECT  2.730 3.290 3.310 3.690 ;
        RECT  2.980 1.000 4.290 1.240 ;
        RECT  2.240 1.210 3.220 1.450 ;
        RECT  1.510 1.340 2.480 1.580 ;
        RECT  1.510 1.260 1.910 1.660 ;
        RECT  1.680 1.340 1.920 4.470 ;
        RECT  1.460 4.070 1.920 4.470 ;
        RECT  4.130 1.560 4.710 1.800 ;
        RECT  4.130 1.560 4.370 2.750 ;
        RECT  4.030 2.510 4.270 3.600 ;
        RECT  4.030 3.350 4.610 3.600 ;
        RECT  3.650 1.480 3.890 2.090 ;
        RECT  5.210 2.530 5.610 2.930 ;
        RECT  4.850 2.860 5.450 3.100 ;
        RECT  3.550 1.850 3.790 4.110 ;
        RECT  4.850 2.860 5.090 4.110 ;
        RECT  3.550 3.870 5.090 4.110 ;
        RECT  4.610 2.050 6.110 2.290 ;
        RECT  4.610 2.050 4.850 2.620 ;
        RECT  5.870 1.510 6.110 3.580 ;
        RECT  5.510 3.340 6.110 3.580 ;
        RECT  7.190 1.100 7.700 1.500 ;
        RECT  7.190 1.100 7.430 3.460 ;
        RECT  7.030 3.060 7.430 3.460 ;
        RECT  6.370 1.460 6.930 1.700 ;
        RECT  7.780 2.610 8.360 2.850 ;
        RECT  6.370 1.460 6.610 3.950 ;
        RECT  7.780 2.610 8.020 3.950 ;
        RECT  6.370 3.710 8.020 3.950 ;
        RECT  7.700 1.910 9.100 2.150 ;
        RECT  8.860 2.330 11.370 2.730 ;
        RECT  8.860 1.300 9.100 3.380 ;
        RECT  8.330 3.140 9.100 3.380 ;
    END
END dfnrq4

MACRO dfnrq2
    CLASS CORE ;
    FOREIGN dfnrq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.145  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.030 3.140 10.580 3.380 ;
        RECT  10.340 1.460 10.580 3.380 ;
        RECT  10.060 1.460 10.580 2.020 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  10.680 4.070 10.920 5.600 ;
        RECT  9.370 4.070 9.610 5.600 ;
        RECT  8.530 4.190 8.770 5.600 ;
        RECT  5.540 4.510 5.780 5.600 ;
        RECT  2.650 4.520 2.890 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  10.650 0.000 11.050 0.890 ;
        RECT  9.290 0.000 9.690 0.890 ;
        RECT  8.090 0.000 8.490 0.890 ;
        RECT  5.490 0.000 5.910 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.700 ;
        RECT  1.590 3.460 2.440 3.700 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.240 2.190 3.480 3.700 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 4.550 4.270 ;
        RECT  4.510 1.660 4.750 3.730 ;
        RECT  4.510 3.330 5.040 3.730 ;
        RECT  3.980 1.180 5.250 1.420 ;
        RECT  3.690 1.600 4.220 2.000 ;
        RECT  5.010 1.180 5.250 3.090 ;
        RECT  5.010 2.850 6.070 3.090 ;
        RECT  3.980 1.180 4.220 3.640 ;
        RECT  5.890 1.770 6.130 2.610 ;
        RECT  5.890 2.370 6.550 2.610 ;
        RECT  6.310 2.370 6.550 4.270 ;
        RECT  4.830 4.030 6.550 4.270 ;
        RECT  7.290 1.690 8.030 1.930 ;
        RECT  7.790 1.690 8.030 4.490 ;
        RECT  8.720 1.100 9.120 1.370 ;
        RECT  6.550 1.130 9.120 1.370 ;
        RECT  6.550 1.130 7.050 2.000 ;
        RECT  6.810 1.130 7.050 2.410 ;
        RECT  7.050 2.170 7.290 4.310 ;
        RECT  8.780 1.610 9.020 2.850 ;
        RECT  8.270 2.430 9.020 2.670 ;
        RECT  8.580 2.610 9.910 2.850 ;
        RECT  8.580 2.430 8.820 3.460 ;
    END
END dfnrq2

MACRO dfnrq1
    CLASS CORE ;
    FOREIGN dfnrq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.076  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.580 3.140 10.490 3.580 ;
        RECT  10.140 1.460 10.490 3.580 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  9.480 4.070 9.720 5.600 ;
        RECT  8.530 4.190 8.770 5.600 ;
        RECT  5.540 4.510 5.780 5.600 ;
        RECT  2.650 4.520 2.890 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  9.320 0.000 9.720 0.890 ;
        RECT  8.090 0.000 8.490 0.890 ;
        RECT  5.490 0.000 5.910 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.700 ;
        RECT  1.590 3.460 2.440 3.700 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.240 2.190 3.480 3.700 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 4.550 4.270 ;
        RECT  4.510 1.660 4.750 3.730 ;
        RECT  4.510 3.330 5.040 3.730 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  3.900 1.180 4.220 2.000 ;
        RECT  3.690 1.600 4.220 2.000 ;
        RECT  5.010 1.180 5.250 3.090 ;
        RECT  5.010 2.850 6.070 3.090 ;
        RECT  3.980 1.180 4.220 3.640 ;
        RECT  5.890 1.770 6.130 2.610 ;
        RECT  5.890 2.370 6.550 2.610 ;
        RECT  6.310 2.370 6.550 4.270 ;
        RECT  4.830 4.030 6.550 4.270 ;
        RECT  7.290 1.610 7.770 2.010 ;
        RECT  7.530 1.610 7.770 4.410 ;
        RECT  7.530 4.170 8.110 4.410 ;
        RECT  8.010 2.430 8.930 2.670 ;
        RECT  8.690 1.610 8.930 3.450 ;
        RECT  6.550 1.130 9.420 1.370 ;
        RECT  6.550 1.130 7.050 2.000 ;
        RECT  6.810 1.130 7.050 2.490 ;
        RECT  9.180 1.130 9.420 2.540 ;
        RECT  7.050 2.250 7.290 4.310 ;
    END
END dfnrq1

MACRO dfnrn4
    CLASS CORE ;
    FOREIGN dfnrn4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.310 2.580 8.910 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.280 2.520 0.520 3.250 ;
        RECT  0.120 3.140 0.500 3.580 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.758  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.370 1.590 11.930 1.830 ;
        RECT  10.440 1.640 11.530 1.880 ;
        RECT  9.700 3.790 11.400 4.030 ;
        RECT  10.660 2.580 11.140 3.020 ;
        RECT  10.660 1.640 10.900 4.030 ;
        RECT  10.040 1.590 10.590 1.830 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.320 5.600 ;
        RECT  11.740 4.390 12.140 5.600 ;
        RECT  10.440 4.400 10.840 5.600 ;
        RECT  9.140 4.400 9.540 5.600 ;
        RECT  7.700 4.710 8.100 5.600 ;
        RECT  5.590 4.710 5.990 5.600 ;
        RECT  2.840 4.710 3.240 5.600 ;
        RECT  0.160 4.080 0.560 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.320 0.740 ;
        RECT  10.790 0.000 11.190 1.370 ;
        RECT  9.300 0.000 9.700 1.370 ;
        RECT  7.820 0.000 8.220 1.420 ;
        RECT  5.830 0.000 6.230 0.890 ;
        RECT  2.960 0.000 3.360 1.750 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 1.220 1.060 2.110 ;
        RECT  0.800 1.880 1.040 3.710 ;
        RECT  2.290 1.240 2.550 1.800 ;
        RECT  2.040 1.560 2.550 1.800 ;
        RECT  2.040 1.560 2.280 2.380 ;
        RECT  2.020 2.180 2.260 3.740 ;
        RECT  2.020 3.500 2.600 3.740 ;
        RECT  1.560 1.200 1.800 2.020 ;
        RECT  3.210 2.520 3.450 3.350 ;
        RECT  2.840 3.110 3.450 3.350 ;
        RECT  1.540 1.910 1.780 4.310 ;
        RECT  2.840 3.110 3.080 4.310 ;
        RECT  1.540 4.060 3.080 4.310 ;
        RECT  3.780 1.620 4.020 2.280 ;
        RECT  2.520 2.040 4.020 2.280 ;
        RECT  2.520 2.040 2.760 2.730 ;
        RECT  3.690 2.040 3.930 4.090 ;
        RECT  3.500 3.690 3.930 4.090 ;
        RECT  4.930 1.990 5.500 2.230 ;
        RECT  5.260 1.610 5.500 2.230 ;
        RECT  4.770 2.000 5.010 3.510 ;
        RECT  4.770 3.270 5.360 3.510 ;
        RECT  4.290 1.520 4.840 1.760 ;
        RECT  5.980 2.960 6.460 3.200 ;
        RECT  6.220 2.500 6.460 3.200 ;
        RECT  5.600 3.120 6.220 3.360 ;
        RECT  4.290 1.520 4.530 3.990 ;
        RECT  5.600 3.120 5.840 3.990 ;
        RECT  4.290 3.750 5.840 3.990 ;
        RECT  5.740 1.610 6.870 1.850 ;
        RECT  6.540 1.680 6.940 2.170 ;
        RECT  5.740 1.610 5.980 2.720 ;
        RECT  5.290 2.470 5.980 2.720 ;
        RECT  5.290 2.470 5.690 2.870 ;
        RECT  6.700 1.680 6.940 3.640 ;
        RECT  6.580 3.430 6.820 3.940 ;
        RECT  6.270 3.700 6.820 3.940 ;
        RECT  4.190 0.980 5.580 1.220 ;
        RECT  6.480 1.020 7.480 1.340 ;
        RECT  5.350 1.130 6.720 1.370 ;
        RECT  7.080 1.020 7.480 1.420 ;
        RECT  7.210 1.020 7.450 3.380 ;
        RECT  7.180 3.170 7.430 3.750 ;
        RECT  8.640 1.290 8.880 2.000 ;
        RECT  7.730 1.760 8.880 2.000 ;
        RECT  7.730 1.760 7.970 4.230 ;
        RECT  7.730 3.260 8.820 3.500 ;
        RECT  7.180 3.990 7.990 4.230 ;
        RECT  7.730 3.260 7.990 4.230 ;
        RECT  5.090 4.230 7.420 4.470 ;
        RECT  4.030 4.380 5.320 4.620 ;
    END
END dfnrn4

MACRO dfnrn2
    CLASS CORE ;
    FOREIGN dfnrn2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.510 0.790 2.910 ;
        RECT  0.120 2.020 0.500 2.910 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.060 1.460 10.580 2.020 ;
        RECT  10.060 1.460 10.430 3.450 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  10.680 4.070 10.920 5.600 ;
        RECT  9.370 4.070 9.610 5.600 ;
        RECT  8.530 4.190 8.770 5.600 ;
        RECT  5.540 4.510 5.780 5.600 ;
        RECT  2.650 4.510 2.890 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  10.650 0.000 11.050 0.890 ;
        RECT  9.290 0.000 9.690 0.890 ;
        RECT  8.090 0.000 8.490 0.890 ;
        RECT  5.490 0.000 5.910 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.700 ;
        RECT  1.590 3.460 2.440 3.700 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.240 2.190 3.480 3.700 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.150 1.270 3.390 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 4.550 4.270 ;
        RECT  4.510 1.660 4.750 3.730 ;
        RECT  4.510 3.330 5.040 3.730 ;
        RECT  3.980 1.180 5.250 1.420 ;
        RECT  3.690 1.600 4.220 2.000 ;
        RECT  5.010 1.180 5.250 3.090 ;
        RECT  5.010 2.850 6.070 3.090 ;
        RECT  3.980 1.180 4.220 3.640 ;
        RECT  5.890 1.770 6.130 2.610 ;
        RECT  5.890 2.370 6.550 2.610 ;
        RECT  6.310 2.370 6.550 4.270 ;
        RECT  4.830 4.030 6.550 4.270 ;
        RECT  7.290 1.690 8.030 1.930 ;
        RECT  7.790 1.690 8.030 4.490 ;
        RECT  8.780 1.610 9.020 2.670 ;
        RECT  8.270 2.430 9.020 2.670 ;
        RECT  8.580 2.430 8.820 3.450 ;
        RECT  6.630 1.130 9.510 1.370 ;
        RECT  6.630 1.130 6.870 2.140 ;
        RECT  6.810 1.900 7.050 2.410 ;
        RECT  9.270 1.130 9.510 2.540 ;
        RECT  7.050 2.170 7.290 4.310 ;
    END
END dfnrn2

MACRO dfnrn1
    CLASS CORE ;
    FOREIGN dfnrn1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.510 0.790 2.910 ;
        RECT  0.120 2.020 0.500 2.910 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.076  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.580 3.140 10.370 3.580 ;
        RECT  9.970 1.460 10.370 3.580 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  9.480 4.070 9.720 5.600 ;
        RECT  8.530 4.190 8.770 5.600 ;
        RECT  5.540 4.510 5.780 5.600 ;
        RECT  2.650 4.510 2.890 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  9.200 0.000 9.600 0.890 ;
        RECT  8.090 0.000 8.490 0.890 ;
        RECT  5.490 0.000 5.910 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.700 ;
        RECT  1.590 3.460 2.440 3.700 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.240 2.190 3.480 3.700 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.150 1.270 3.390 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 4.550 4.270 ;
        RECT  4.510 1.660 4.750 3.730 ;
        RECT  4.510 3.330 5.040 3.730 ;
        RECT  3.980 1.180 5.250 1.420 ;
        RECT  3.690 1.600 4.220 2.000 ;
        RECT  5.010 1.180 5.250 3.090 ;
        RECT  5.010 2.850 6.070 3.090 ;
        RECT  3.980 1.180 4.220 3.640 ;
        RECT  5.890 1.770 6.130 2.610 ;
        RECT  5.890 2.370 6.550 2.610 ;
        RECT  6.310 2.370 6.550 4.270 ;
        RECT  4.830 4.030 6.550 4.270 ;
        RECT  7.290 1.610 7.770 2.010 ;
        RECT  7.530 1.610 7.770 4.410 ;
        RECT  7.530 4.170 8.110 4.410 ;
        RECT  8.010 2.430 8.930 2.670 ;
        RECT  8.690 1.610 8.930 3.450 ;
        RECT  6.550 1.130 9.420 1.370 ;
        RECT  6.550 1.130 7.050 2.000 ;
        RECT  6.790 1.130 7.050 2.490 ;
        RECT  9.180 1.130 9.420 2.540 ;
        RECT  7.050 2.250 7.290 4.310 ;
    END
END dfnrn1

MACRO dfnrb4
    CLASS CORE ;
    FOREIGN dfnrb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.390 2.340 0.790 2.740 ;
        RECT  0.120 2.580 0.640 2.820 ;
        RECT  0.120 2.580 0.500 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.770 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.807  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.420 1.290 11.300 1.690 ;
        RECT  10.900 1.120 11.300 1.690 ;
        RECT  9.390 2.820 11.140 3.220 ;
        RECT  10.700 2.580 11.140 3.220 ;
        RECT  10.740 1.290 11.140 3.220 ;
        RECT  9.420 1.070 9.820 1.690 ;
        RECT  9.390 2.820 9.790 4.620 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.235  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.860 1.050 14.260 1.740 ;
        RECT  13.540 1.500 13.940 3.020 ;
        RECT  13.150 2.580 13.550 3.720 ;
        RECT  12.380 1.500 13.940 1.900 ;
        RECT  11.850 2.580 13.940 2.980 ;
        RECT  12.380 1.050 12.780 1.900 ;
        RECT  11.850 2.580 12.250 3.780 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 14.560 5.600 ;
        RECT  13.930 4.090 14.330 5.600 ;
        RECT  12.590 4.170 12.990 5.600 ;
        RECT  11.290 4.170 11.690 5.600 ;
        RECT  10.030 3.520 10.270 5.600 ;
        RECT  8.650 4.330 9.050 5.600 ;
        RECT  7.380 4.300 7.780 5.600 ;
        RECT  4.640 4.710 5.040 5.600 ;
        RECT  1.990 4.220 2.390 5.600 ;
        RECT  0.720 4.150 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 14.560 0.740 ;
        RECT  13.120 0.000 13.520 0.980 ;
        RECT  11.640 0.000 12.040 0.980 ;
        RECT  10.160 0.000 10.560 0.980 ;
        RECT  7.980 0.000 8.380 1.730 ;
        RECT  5.020 0.000 5.420 1.640 ;
        RECT  2.170 0.000 2.570 0.890 ;
        RECT  0.920 0.000 1.320 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.820 1.290 2.060 ;
        RECT  1.050 2.520 1.480 2.920 ;
        RECT  1.050 1.820 1.290 3.140 ;
        RECT  0.970 2.900 1.210 3.500 ;
        RECT  0.150 3.260 1.210 3.500 ;
        RECT  2.780 1.630 3.280 2.030 ;
        RECT  3.040 1.630 3.280 3.790 ;
        RECT  2.730 3.550 3.280 3.790 ;
        RECT  3.050 0.980 4.300 1.220 ;
        RECT  1.590 1.130 3.290 1.370 ;
        RECT  1.590 1.130 1.830 2.300 ;
        RECT  1.720 2.060 1.960 3.920 ;
        RECT  1.460 3.520 1.960 3.920 ;
        RECT  4.080 1.700 4.680 1.940 ;
        RECT  4.080 1.700 4.320 2.490 ;
        RECT  4.050 2.250 4.310 3.870 ;
        RECT  4.050 3.470 4.450 3.870 ;
        RECT  3.600 1.570 3.840 2.120 ;
        RECT  5.400 2.450 5.640 3.360 ;
        RECT  4.770 3.120 5.640 3.360 ;
        RECT  3.570 1.990 3.810 4.350 ;
        RECT  4.770 3.120 5.010 4.350 ;
        RECT  3.290 4.110 5.010 4.350 ;
        RECT  3.290 4.110 3.690 4.620 ;
        RECT  4.920 1.970 6.080 2.210 ;
        RECT  5.840 1.480 6.080 2.210 ;
        RECT  4.920 1.970 5.160 2.540 ;
        RECT  4.560 2.300 5.160 2.540 ;
        RECT  4.560 2.300 4.800 2.850 ;
        RECT  5.880 1.980 6.120 3.960 ;
        RECT  5.410 3.720 6.120 3.960 ;
        RECT  7.060 1.590 7.640 1.830 ;
        RECT  7.060 1.590 7.300 2.550 ;
        RECT  6.860 2.310 7.100 3.320 ;
        RECT  6.580 1.510 6.820 2.070 ;
        RECT  8.320 2.450 8.560 3.180 ;
        RECT  7.340 2.940 8.560 3.180 ;
        RECT  7.340 2.940 7.580 3.800 ;
        RECT  6.360 3.560 7.580 3.800 ;
        RECT  6.360 1.830 6.600 4.620 ;
        RECT  6.010 4.380 6.600 4.620 ;
        RECT  7.840 1.970 10.500 2.210 ;
        RECT  8.800 1.930 10.500 2.330 ;
        RECT  7.540 2.090 8.080 2.490 ;
        RECT  8.800 1.560 9.040 3.660 ;
        RECT  8.120 3.420 9.040 3.660 ;
    END
END dfnrb4

MACRO dfnrb2
    CLASS CORE ;
    FOREIGN dfnrb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.440 0.790 2.840 ;
        RECT  0.120 2.020 0.500 2.840 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.318  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.330 3.330 11.140 3.580 ;
        RECT  10.700 3.140 11.140 3.580 ;
        RECT  10.700 1.620 10.940 3.580 ;
        RECT  10.300 1.620 10.940 1.860 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.189  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.760 3.330 12.760 3.570 ;
        RECT  12.370 1.850 12.760 3.570 ;
        RECT  11.760 1.850 12.760 2.090 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.880 5.600 ;
        RECT  12.410 4.280 12.650 5.600 ;
        RECT  11.100 4.290 11.340 5.600 ;
        RECT  9.790 4.290 10.030 5.600 ;
        RECT  8.760 4.400 9.000 5.600 ;
        RECT  5.540 4.510 5.780 5.600 ;
        RECT  2.650 4.510 2.890 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.880 0.740 ;
        RECT  12.330 0.000 12.730 0.890 ;
        RECT  10.970 0.000 11.370 0.890 ;
        RECT  9.610 0.000 10.010 0.890 ;
        RECT  8.140 0.000 8.540 0.890 ;
        RECT  5.490 0.000 5.910 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.700 ;
        RECT  1.590 3.460 2.440 3.700 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.240 2.190 3.480 3.700 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 4.550 4.270 ;
        RECT  4.510 1.660 4.750 3.730 ;
        RECT  4.510 3.330 5.040 3.730 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  3.900 1.180 4.220 2.000 ;
        RECT  3.690 1.600 4.220 2.000 ;
        RECT  5.010 1.180 5.250 3.090 ;
        RECT  5.010 2.850 6.070 3.090 ;
        RECT  3.980 1.180 4.220 3.640 ;
        RECT  5.890 1.770 6.130 2.610 ;
        RECT  5.890 2.370 6.550 2.610 ;
        RECT  6.310 2.370 6.550 4.270 ;
        RECT  4.830 4.030 6.550 4.270 ;
        RECT  7.290 1.610 7.660 2.010 ;
        RECT  7.420 1.610 7.660 4.620 ;
        RECT  7.420 4.380 7.970 4.620 ;
        RECT  8.990 1.610 9.230 3.040 ;
        RECT  8.060 2.590 9.230 2.830 ;
        RECT  8.730 2.800 10.430 3.040 ;
        RECT  8.730 2.590 8.970 3.450 ;
        RECT  8.700 1.080 9.070 1.370 ;
        RECT  6.550 1.130 11.500 1.370 ;
        RECT  6.550 1.130 7.050 2.000 ;
        RECT  11.260 1.130 11.500 2.710 ;
        RECT  6.810 1.130 7.050 2.490 ;
        RECT  11.260 2.470 11.910 2.710 ;
        RECT  6.910 2.250 7.150 4.620 ;
    END
END dfnrb2

MACRO dfnrb1
    CLASS CORE ;
    FOREIGN dfnrb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.440 0.790 2.840 ;
        RECT  0.120 2.020 0.500 2.840 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.000  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.430 2.020 10.050 2.460 ;
        RECT  9.430 1.610 9.670 3.450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.016  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.140 3.140 11.050 3.580 ;
        RECT  10.650 1.540 11.050 3.580 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  10.160 4.070 10.400 5.600 ;
        RECT  8.500 4.400 8.740 5.600 ;
        RECT  5.540 4.510 5.780 5.600 ;
        RECT  2.650 4.510 2.890 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  10.050 0.000 10.450 0.890 ;
        RECT  7.880 0.000 8.280 0.890 ;
        RECT  5.490 0.000 5.910 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.700 ;
        RECT  1.590 3.460 2.440 3.700 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.240 2.190 3.480 3.700 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 4.550 4.270 ;
        RECT  4.510 1.660 4.750 3.730 ;
        RECT  4.510 3.330 5.040 3.730 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  3.900 1.180 4.220 2.000 ;
        RECT  3.690 1.600 4.220 2.000 ;
        RECT  5.010 1.180 5.250 3.090 ;
        RECT  5.010 2.850 6.070 3.090 ;
        RECT  3.980 1.180 4.220 3.640 ;
        RECT  5.890 1.770 6.130 2.610 ;
        RECT  5.890 2.370 6.550 2.610 ;
        RECT  6.310 2.370 6.550 4.270 ;
        RECT  4.830 4.030 6.550 4.270 ;
        RECT  7.290 1.610 7.660 2.010 ;
        RECT  7.420 1.610 7.660 4.620 ;
        RECT  7.420 4.380 7.970 4.620 ;
        RECT  8.440 1.080 8.810 1.370 ;
        RECT  6.550 1.130 8.810 1.370 ;
        RECT  6.550 1.130 7.050 2.000 ;
        RECT  6.810 1.130 7.050 2.490 ;
        RECT  6.910 2.250 7.150 4.620 ;
        RECT  8.730 1.610 8.970 2.830 ;
        RECT  8.010 2.590 8.970 2.830 ;
        RECT  8.560 2.590 8.800 3.450 ;
    END
END dfnrb1

MACRO dfnfb4
    CLASS CORE ;
    FOREIGN dfnfb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.360 2.360 0.800 2.770 ;
        RECT  0.120 2.530 0.580 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.380  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.360 2.740 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.838  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.260 2.020 11.730 2.460 ;
        RECT  9.720 2.990 11.650 3.230 ;
        RECT  11.410 1.610 11.650 3.230 ;
        RECT  11.260 1.610 11.650 2.460 ;
        RECT  11.020 2.990 11.260 4.320 ;
        RECT  9.190 1.610 11.650 1.850 ;
        RECT  10.570 1.290 10.810 1.850 ;
        RECT  9.720 2.990 9.960 4.320 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.833  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.870 2.450 14.110 3.550 ;
        RECT  12.080 2.450 14.110 2.690 ;
        RECT  12.940 2.020 13.800 2.690 ;
        RECT  13.560 1.110 13.800 2.690 ;
        RECT  12.390 2.450 12.630 4.320 ;
        RECT  12.080 0.980 12.320 2.690 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.120 5.600 ;
        RECT  14.540 4.150 14.940 5.600 ;
        RECT  13.060 4.050 13.420 5.600 ;
        RECT  11.690 4.610 12.090 5.600 ;
        RECT  10.380 4.610 10.780 5.600 ;
        RECT  9.070 4.610 9.470 5.600 ;
        RECT  7.630 4.420 8.030 5.600 ;
        RECT  4.940 4.290 5.340 5.600 ;
        RECT  2.140 4.710 2.540 5.600 ;
        RECT  0.720 4.090 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.120 0.740 ;
        RECT  12.740 0.000 13.140 0.980 ;
        RECT  11.260 0.000 11.660 1.200 ;
        RECT  9.790 0.000 10.190 0.890 ;
        RECT  7.460 0.000 7.860 1.110 ;
        RECT  4.610 0.000 5.010 0.890 ;
        RECT  2.340 0.000 2.740 1.090 ;
        RECT  0.880 0.000 1.280 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.140 1.840 1.280 2.080 ;
        RECT  1.040 1.840 1.280 2.920 ;
        RECT  1.040 2.520 1.500 2.920 ;
        RECT  1.160 2.520 1.400 3.500 ;
        RECT  0.150 3.260 1.400 3.500 ;
        RECT  2.810 1.460 3.220 1.860 ;
        RECT  2.980 1.460 3.220 3.660 ;
        RECT  2.740 3.260 3.220 3.660 ;
        RECT  4.110 1.610 4.690 1.850 ;
        RECT  4.110 1.610 4.350 2.590 ;
        RECT  4.160 2.350 4.400 3.450 ;
        RECT  5.250 0.980 5.810 1.220 ;
        RECT  3.630 1.130 5.490 1.370 ;
        RECT  3.630 1.130 3.870 2.340 ;
        RECT  3.560 2.100 3.800 4.140 ;
        RECT  5.580 1.670 6.050 2.070 ;
        RECT  4.640 2.300 4.880 3.080 ;
        RECT  4.640 2.840 5.820 3.080 ;
        RECT  5.580 1.670 5.820 3.450 ;
        RECT  1.520 1.000 2.090 1.240 ;
        RECT  1.520 1.000 1.770 2.070 ;
        RECT  4.240 3.810 5.950 4.050 ;
        RECT  1.740 1.670 1.980 4.470 ;
        RECT  1.460 4.070 1.980 4.470 ;
        RECT  5.710 3.810 5.950 4.620 ;
        RECT  1.460 4.230 3.170 4.470 ;
        RECT  4.240 3.810 4.480 4.620 ;
        RECT  2.930 4.380 4.480 4.620 ;
        RECT  5.710 4.380 6.450 4.620 ;
        RECT  6.970 1.570 7.530 1.810 ;
        RECT  6.970 1.570 7.210 3.450 ;
        RECT  6.970 3.050 7.430 3.450 ;
        RECT  6.470 1.610 6.710 2.320 ;
        RECT  8.140 2.520 8.380 3.480 ;
        RECT  7.670 3.240 8.380 3.480 ;
        RECT  6.370 2.080 6.610 4.140 ;
        RECT  7.670 3.240 7.910 4.140 ;
        RECT  6.370 3.900 7.910 4.140 ;
        RECT  7.770 1.710 8.890 1.950 ;
        RECT  8.490 1.630 8.890 2.030 ;
        RECT  8.650 1.630 8.890 2.660 ;
        RECT  7.770 1.710 8.010 2.290 ;
        RECT  7.460 2.050 8.010 2.290 ;
        RECT  8.650 2.260 10.880 2.660 ;
        RECT  7.460 2.050 7.700 2.700 ;
        RECT  9.220 2.260 9.460 4.060 ;
        RECT  8.370 3.820 9.460 4.060 ;
    END
END dfnfb4

MACRO dfnfb2
    CLASS CORE ;
    FOREIGN dfnfb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.070 2.660 1.650 3.030 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.370 2.580 2.720 3.190 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.318  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.330 3.330 11.140 3.580 ;
        RECT  10.700 3.140 11.140 3.580 ;
        RECT  10.700 1.620 10.940 3.580 ;
        RECT  10.300 1.620 10.940 1.860 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.189  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.760 3.330 12.760 3.570 ;
        RECT  12.370 1.850 12.760 3.570 ;
        RECT  11.760 1.850 12.760 2.090 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.880 5.600 ;
        RECT  12.410 4.280 12.650 5.600 ;
        RECT  11.100 4.290 11.340 5.600 ;
        RECT  9.790 4.290 10.030 5.600 ;
        RECT  8.760 4.400 9.000 5.600 ;
        RECT  5.540 4.340 5.780 5.600 ;
        RECT  2.650 4.420 2.890 5.600 ;
        RECT  0.550 4.150 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.880 0.740 ;
        RECT  12.330 0.000 12.730 0.890 ;
        RECT  10.970 0.000 11.370 0.890 ;
        RECT  9.610 0.000 10.010 0.890 ;
        RECT  8.140 0.000 8.540 0.890 ;
        RECT  5.490 0.000 5.910 1.260 ;
        RECT  2.210 1.680 2.770 1.920 ;
        RECT  2.530 0.000 2.770 1.920 ;
        RECT  0.720 0.000 1.120 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.290 1.220 ;
        RECT  1.590 0.980 1.830 2.420 ;
        RECT  0.660 1.940 1.830 2.180 ;
        RECT  1.590 2.150 2.130 2.420 ;
        RECT  0.660 1.940 0.900 2.490 ;
        RECT  1.890 2.150 2.130 3.700 ;
        RECT  1.510 3.460 2.440 3.700 ;
        RECT  3.030 1.660 3.270 2.530 ;
        RECT  3.240 2.290 3.480 3.700 ;
        RECT  0.120 1.320 0.550 1.700 ;
        RECT  0.120 1.320 0.360 3.800 ;
        RECT  0.120 3.400 1.270 3.800 ;
        RECT  1.030 3.400 1.270 4.180 ;
        RECT  1.030 3.940 4.550 4.180 ;
        RECT  4.150 3.940 4.550 4.350 ;
        RECT  4.510 1.660 4.750 3.560 ;
        RECT  4.510 3.320 5.060 3.560 ;
        RECT  3.980 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.810 ;
        RECT  5.010 1.570 5.620 1.810 ;
        RECT  3.690 1.600 4.220 2.000 ;
        RECT  5.380 1.570 5.620 3.090 ;
        RECT  5.380 2.850 6.070 3.090 ;
        RECT  3.980 1.180 4.220 3.640 ;
        RECT  5.890 1.770 6.130 2.610 ;
        RECT  5.890 2.370 6.550 2.610 ;
        RECT  6.310 2.370 6.550 4.100 ;
        RECT  4.830 3.860 6.550 4.100 ;
        RECT  4.830 3.860 5.230 4.350 ;
        RECT  7.290 1.610 7.660 2.010 ;
        RECT  7.420 1.610 7.660 4.620 ;
        RECT  7.420 4.380 7.970 4.620 ;
        RECT  8.990 1.610 9.230 3.040 ;
        RECT  8.060 2.590 9.230 2.830 ;
        RECT  8.730 2.800 10.430 3.040 ;
        RECT  8.730 2.590 8.970 3.450 ;
        RECT  8.700 1.080 9.070 1.370 ;
        RECT  6.630 1.130 11.500 1.370 ;
        RECT  6.630 1.130 6.870 2.140 ;
        RECT  11.260 1.130 11.500 2.710 ;
        RECT  6.810 1.900 7.050 2.490 ;
        RECT  11.260 2.470 11.910 2.710 ;
        RECT  6.910 2.250 7.150 4.620 ;
    END
END dfnfb2

MACRO dfnfb1
    CLASS CORE ;
    FOREIGN dfnfb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.070 2.660 1.650 3.030 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.370 2.580 2.720 3.190 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.009  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.430 2.020 10.050 2.460 ;
        RECT  9.430 1.610 9.670 3.450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.991  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.140 3.140 11.050 3.580 ;
        RECT  10.650 1.590 11.050 3.580 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  10.160 4.070 10.400 5.600 ;
        RECT  8.500 4.400 8.740 5.600 ;
        RECT  5.540 4.340 5.780 5.600 ;
        RECT  2.650 4.420 2.890 5.600 ;
        RECT  0.550 4.150 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  10.050 0.000 10.450 0.890 ;
        RECT  7.880 0.000 8.280 0.890 ;
        RECT  5.490 0.000 5.910 1.260 ;
        RECT  2.210 1.680 2.770 1.920 ;
        RECT  2.530 0.000 2.770 1.920 ;
        RECT  0.720 0.000 1.120 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.290 1.220 ;
        RECT  1.590 0.980 1.830 2.420 ;
        RECT  0.660 1.940 1.830 2.180 ;
        RECT  1.590 2.150 2.130 2.420 ;
        RECT  0.660 1.940 0.900 2.490 ;
        RECT  1.890 2.150 2.130 3.700 ;
        RECT  1.510 3.460 2.440 3.700 ;
        RECT  3.030 1.660 3.270 2.530 ;
        RECT  3.240 2.290 3.480 3.700 ;
        RECT  0.120 1.320 0.550 1.700 ;
        RECT  0.120 1.320 0.360 3.800 ;
        RECT  0.120 3.400 1.270 3.800 ;
        RECT  1.030 3.400 1.270 4.180 ;
        RECT  1.030 3.940 4.550 4.180 ;
        RECT  4.150 3.940 4.550 4.350 ;
        RECT  4.510 1.660 4.750 3.560 ;
        RECT  4.510 3.320 5.060 3.560 ;
        RECT  3.980 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.810 ;
        RECT  5.010 1.570 5.620 1.810 ;
        RECT  3.690 1.600 4.220 2.000 ;
        RECT  5.380 1.570 5.620 3.090 ;
        RECT  5.380 2.850 6.070 3.090 ;
        RECT  3.980 1.180 4.220 3.640 ;
        RECT  5.890 1.770 6.130 2.610 ;
        RECT  5.890 2.370 6.550 2.610 ;
        RECT  6.310 2.370 6.550 4.100 ;
        RECT  4.830 3.860 6.550 4.100 ;
        RECT  4.830 3.860 5.230 4.350 ;
        RECT  7.290 1.610 7.660 2.010 ;
        RECT  7.420 1.610 7.660 4.620 ;
        RECT  7.420 4.380 7.970 4.620 ;
        RECT  8.440 1.080 8.810 1.370 ;
        RECT  6.630 1.130 8.810 1.370 ;
        RECT  6.630 1.130 6.870 2.140 ;
        RECT  6.810 1.900 7.050 2.490 ;
        RECT  6.910 2.250 7.150 4.620 ;
        RECT  8.730 1.610 8.970 2.830 ;
        RECT  8.010 2.590 8.970 2.830 ;
        RECT  8.560 2.590 8.800 3.450 ;
    END
END dfnfb1

MACRO dfcrq4
    CLASS CORE ;
    FOREIGN dfcrq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 2.520 6.160 3.020 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.440 2.160 0.680 2.770 ;
        RECT  0.120 2.530 0.580 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.360 2.740 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.340 2.690 13.320 2.930 ;
        RECT  12.940 1.470 13.320 2.930 ;
        RECT  12.890 1.470 13.320 1.870 ;
        RECT  11.420 1.550 13.320 1.790 ;
        RECT  12.260 3.890 12.660 4.290 ;
        RECT  12.340 2.690 12.580 4.290 ;
        RECT  10.960 3.970 12.660 4.210 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 13.440 5.600 ;
        RECT  12.940 3.170 13.260 5.600 ;
        RECT  12.860 3.170 13.260 3.570 ;
        RECT  11.700 4.620 12.100 5.600 ;
        RECT  10.390 4.620 10.790 5.600 ;
        RECT  8.760 4.650 9.160 5.600 ;
        RECT  4.690 4.710 5.090 5.600 ;
        RECT  2.140 4.710 2.540 5.600 ;
        RECT  0.720 4.150 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 13.440 0.740 ;
        RECT  12.010 0.000 12.410 0.890 ;
        RECT  10.830 0.000 11.230 0.890 ;
        RECT  8.820 0.000 9.220 1.090 ;
        RECT  4.590 0.000 4.990 0.890 ;
        RECT  1.680 0.000 2.080 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.670 1.160 1.910 ;
        RECT  0.920 1.670 1.160 2.590 ;
        RECT  1.160 2.350 1.400 3.500 ;
        RECT  0.150 3.260 1.400 3.500 ;
        RECT  2.800 1.490 3.220 1.890 ;
        RECT  2.980 1.490 3.220 3.840 ;
        RECT  2.740 3.440 3.220 3.840 ;
        RECT  4.110 1.610 4.680 1.850 ;
        RECT  4.110 1.610 4.350 3.500 ;
        RECT  4.110 3.260 5.970 3.500 ;
        RECT  3.620 1.490 3.860 4.080 ;
        RECT  6.470 1.940 6.710 3.990 ;
        RECT  3.550 3.750 6.710 3.990 ;
        RECT  3.550 3.680 3.950 4.080 ;
        RECT  5.720 1.460 7.210 1.700 ;
        RECT  4.960 1.610 5.960 1.850 ;
        RECT  4.960 1.610 5.200 2.730 ;
        RECT  4.590 2.490 5.200 2.730 ;
        RECT  6.970 1.460 7.210 3.820 ;
        RECT  5.240 0.980 7.650 1.220 ;
        RECT  2.320 1.010 4.350 1.250 ;
        RECT  1.590 1.130 2.560 1.370 ;
        RECT  4.110 1.130 5.480 1.370 ;
        RECT  1.590 1.130 1.830 2.170 ;
        RECT  1.640 2.000 1.880 4.470 ;
        RECT  1.460 4.060 1.880 4.470 ;
        RECT  1.460 4.230 3.170 4.470 ;
        RECT  4.200 4.230 7.370 4.470 ;
        RECT  2.930 4.380 4.440 4.620 ;
        RECT  7.130 4.380 8.290 4.620 ;
        RECT  8.310 1.490 8.550 3.450 ;
        RECT  8.310 3.050 8.790 3.450 ;
        RECT  7.480 1.550 7.960 1.950 ;
        RECT  9.490 1.990 9.730 3.480 ;
        RECT  9.140 3.240 9.730 3.480 ;
        RECT  7.720 1.550 7.960 4.140 ;
        RECT  9.140 3.240 9.380 4.140 ;
        RECT  7.720 3.900 9.380 4.140 ;
        RECT  8.810 1.510 10.310 1.750 ;
        RECT  8.810 1.510 9.050 2.540 ;
        RECT  10.070 2.200 12.060 2.600 ;
        RECT  10.070 1.510 10.310 4.240 ;
        RECT  9.620 4.000 10.310 4.240 ;
    END
END dfcrq4

MACRO dfcrq2
    CLASS CORE ;
    FOREIGN dfcrq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.020 5.460 2.770 ;
        RECT  5.000 2.500 5.240 3.160 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.791  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.230 1.770 12.170 2.170 ;
        RECT  10.700 3.770 12.090 4.010 ;
        RECT  11.850 1.770 12.090 4.010 ;
        RECT  10.700 3.700 11.140 4.140 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.320 5.600 ;
        RECT  11.770 4.610 12.170 5.600 ;
        RECT  10.540 4.380 10.780 5.600 ;
        RECT  9.170 4.510 9.410 5.600 ;
        RECT  6.450 4.710 6.850 5.600 ;
        RECT  5.260 4.710 5.660 5.600 ;
        RECT  2.340 4.710 2.740 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.320 0.740 ;
        RECT  10.610 0.000 11.550 0.980 ;
        RECT  8.880 0.000 9.280 0.980 ;
        RECT  5.940 0.000 6.180 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.710 ;
        RECT  1.590 3.470 2.430 3.710 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.230 2.190 3.470 3.730 ;
        RECT  4.510 1.660 4.750 3.720 ;
        RECT  5.480 3.220 6.370 3.460 ;
        RECT  4.510 3.400 5.720 3.720 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.740 ;
        RECT  5.010 1.500 6.420 1.740 ;
        RECT  3.900 1.180 4.210 2.000 ;
        RECT  3.690 1.600 4.210 2.000 ;
        RECT  6.180 1.500 6.420 2.500 ;
        RECT  6.180 2.260 6.730 2.500 ;
        RECT  3.970 1.180 4.210 3.730 ;
        RECT  6.710 1.470 6.950 2.020 ;
        RECT  6.710 1.780 7.210 2.020 ;
        RECT  5.700 2.420 5.940 2.980 ;
        RECT  6.970 1.780 7.210 2.980 ;
        RECT  5.700 2.740 7.400 2.980 ;
        RECT  7.160 2.740 7.400 3.730 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 2.390 4.270 ;
        RECT  2.150 4.220 7.270 4.460 ;
        RECT  7.050 4.320 7.980 4.560 ;
        RECT  8.110 1.770 8.720 2.010 ;
        RECT  8.480 1.770 8.720 2.660 ;
        RECT  8.380 2.420 8.620 4.030 ;
        RECT  8.380 3.790 8.960 4.030 ;
        RECT  7.450 1.290 9.380 1.530 ;
        RECT  7.450 1.290 7.690 2.490 ;
        RECT  9.130 1.290 9.380 2.490 ;
        RECT  7.450 2.250 8.140 2.490 ;
        RECT  9.130 2.250 10.300 2.490 ;
        RECT  10.060 2.250 10.300 2.820 ;
        RECT  7.900 2.250 8.140 4.000 ;
        RECT  9.910 1.690 10.780 1.930 ;
        RECT  10.540 1.690 10.780 2.620 ;
        RECT  10.540 2.380 11.050 2.620 ;
        RECT  8.860 3.050 9.920 3.300 ;
        RECT  10.810 2.380 11.050 3.300 ;
        RECT  8.860 3.060 11.050 3.300 ;
        RECT  9.980 3.060 10.220 3.900 ;
    END
END dfcrq2

MACRO dfcrq1
    CLASS CORE ;
    FOREIGN dfcrq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.020 5.460 2.770 ;
        RECT  5.000 2.500 5.240 3.160 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.031  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.700 3.610 11.610 4.140 ;
        RECT  11.290 1.210 11.530 4.140 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.760 5.600 ;
        RECT  10.720 4.380 10.960 5.600 ;
        RECT  9.420 3.530 9.660 5.600 ;
        RECT  6.450 4.710 6.850 5.600 ;
        RECT  5.260 4.710 5.660 5.600 ;
        RECT  2.350 4.710 2.750 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.760 0.740 ;
        RECT  10.610 0.000 11.010 0.980 ;
        RECT  8.880 0.000 9.280 0.980 ;
        RECT  5.940 0.000 6.180 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.710 ;
        RECT  1.590 3.470 2.430 3.710 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.230 2.190 3.470 3.730 ;
        RECT  4.510 1.660 4.750 3.720 ;
        RECT  5.480 3.220 6.370 3.460 ;
        RECT  4.510 3.400 5.720 3.720 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.740 ;
        RECT  5.010 1.500 6.420 1.740 ;
        RECT  3.900 1.180 4.210 2.000 ;
        RECT  3.690 1.600 4.210 2.000 ;
        RECT  6.180 1.500 6.420 2.500 ;
        RECT  6.180 2.260 6.730 2.500 ;
        RECT  3.970 1.180 4.210 3.730 ;
        RECT  6.710 1.470 6.950 2.020 ;
        RECT  6.710 1.780 7.210 2.020 ;
        RECT  5.700 2.420 5.940 2.980 ;
        RECT  6.970 1.780 7.210 2.980 ;
        RECT  5.700 2.740 7.400 2.980 ;
        RECT  7.160 2.740 7.400 3.730 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 2.390 4.270 ;
        RECT  2.150 4.220 7.270 4.460 ;
        RECT  7.050 4.320 7.980 4.560 ;
        RECT  8.110 1.770 8.720 2.010 ;
        RECT  8.480 1.770 8.720 2.660 ;
        RECT  8.380 2.420 8.620 4.030 ;
        RECT  8.380 3.790 8.960 4.030 ;
        RECT  7.450 1.290 9.380 1.530 ;
        RECT  7.450 1.290 7.690 2.490 ;
        RECT  9.130 1.290 9.380 2.490 ;
        RECT  7.450 2.250 8.140 2.490 ;
        RECT  9.130 2.250 10.540 2.490 ;
        RECT  10.300 2.250 10.540 2.820 ;
        RECT  7.900 2.250 8.140 4.000 ;
        RECT  9.910 1.550 11.050 1.790 ;
        RECT  9.910 1.550 10.310 2.010 ;
        RECT  8.860 3.050 10.220 3.290 ;
        RECT  10.810 1.550 11.050 3.300 ;
        RECT  9.980 3.060 11.050 3.300 ;
        RECT  9.980 3.050 10.220 4.620 ;
    END
END dfcrq1

MACRO dfcrn4
    CLASS CORE ;
    FOREIGN dfcrn4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.888  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.250 1.130 9.490 2.940 ;
        RECT  8.700 1.130 9.490 1.370 ;
        RECT  6.190 1.100 8.860 1.340 ;
        RECT  5.300 1.130 6.430 1.370 ;
        RECT  5.100 1.460 5.540 1.900 ;
        RECT  5.300 1.130 5.540 1.900 ;
        RECT  5.270 1.460 5.510 2.860 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.500 0.620 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 2.020 2.740 2.460 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.213  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.740 1.680 12.620 1.920 ;
        RECT  12.320 2.820 12.560 4.430 ;
        RECT  10.950 2.820 12.560 3.060 ;
        RECT  11.820 1.680 12.260 3.060 ;
        RECT  10.950 2.820 11.190 4.350 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 13.440 5.600 ;
        RECT  12.890 4.620 13.290 5.600 ;
        RECT  11.470 3.300 11.870 5.600 ;
        RECT  10.300 4.620 10.700 5.600 ;
        RECT  8.900 4.530 9.300 5.600 ;
        RECT  6.020 4.610 6.420 5.600 ;
        RECT  4.720 4.620 5.120 5.600 ;
        RECT  2.090 4.290 2.490 5.600 ;
        RECT  0.720 4.380 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 13.440 0.740 ;
        RECT  11.480 0.000 11.880 1.170 ;
        RECT  8.980 0.000 9.380 0.890 ;
        RECT  5.510 0.000 5.930 0.890 ;
        RECT  1.720 0.000 2.120 0.890 ;
        RECT  0.920 0.000 1.320 0.900 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.490 1.210 1.730 ;
        RECT  0.970 2.150 1.500 2.550 ;
        RECT  0.970 1.490 1.210 3.800 ;
        RECT  0.150 3.560 1.210 3.800 ;
        RECT  2.800 1.460 3.220 1.780 ;
        RECT  2.980 1.460 3.220 3.160 ;
        RECT  2.910 2.920 3.150 3.930 ;
        RECT  2.390 0.980 4.170 1.220 ;
        RECT  2.320 1.050 2.630 1.290 ;
        RECT  2.320 1.050 2.560 1.610 ;
        RECT  1.510 1.370 2.560 1.610 ;
        RECT  1.510 1.370 1.980 1.780 ;
        RECT  1.740 2.740 2.130 3.140 ;
        RECT  1.740 1.370 1.980 3.860 ;
        RECT  1.450 3.460 1.980 3.860 ;
        RECT  4.360 1.490 4.600 2.360 ;
        RECT  3.940 2.120 4.600 2.360 ;
        RECT  3.940 2.120 4.180 3.890 ;
        RECT  3.940 3.650 5.890 3.890 ;
        RECT  3.460 1.460 3.940 1.850 ;
        RECT  6.230 2.770 6.470 3.780 ;
        RECT  3.460 1.460 3.700 4.620 ;
        RECT  6.150 3.540 6.390 4.370 ;
        RECT  3.460 4.130 6.390 4.370 ;
        RECT  3.390 4.220 3.800 4.620 ;
        RECT  6.180 1.670 6.420 2.530 ;
        RECT  5.750 2.290 6.950 2.530 ;
        RECT  4.420 2.820 4.660 3.410 ;
        RECT  5.650 3.060 5.990 3.300 ;
        RECT  5.750 2.290 5.990 3.300 ;
        RECT  4.420 3.170 5.860 3.410 ;
        RECT  6.710 2.290 6.950 4.090 ;
        RECT  6.870 3.860 7.110 4.410 ;
        RECT  8.470 1.610 8.710 2.350 ;
        RECT  7.670 2.110 8.710 2.350 ;
        RECT  7.670 1.580 7.910 2.950 ;
        RECT  7.670 2.710 8.210 2.950 ;
        RECT  7.970 2.710 8.210 3.810 ;
        RECT  7.970 3.570 8.530 3.810 ;
        RECT  9.730 1.000 10.610 1.240 ;
        RECT  8.530 2.610 8.770 3.330 ;
        RECT  8.770 3.090 9.010 3.810 ;
        RECT  9.470 3.410 9.980 3.810 ;
        RECT  9.730 1.000 9.980 3.810 ;
        RECT  8.770 3.570 9.980 3.810 ;
        RECT  6.840 1.660 7.430 1.900 ;
        RECT  10.220 2.180 11.160 2.580 ;
        RECT  7.190 1.660 7.430 3.430 ;
        RECT  7.190 3.190 7.710 3.430 ;
        RECT  7.470 3.190 7.710 4.290 ;
        RECT  10.220 2.180 10.460 4.290 ;
        RECT  7.470 4.050 10.460 4.290 ;
    END
END dfcrn4

MACRO dfcrn2
    CLASS CORE ;
    FOREIGN dfcrn2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.020 5.460 2.770 ;
        RECT  5.000 2.500 5.240 3.160 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.791  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.230 1.770 12.170 2.170 ;
        RECT  10.700 3.770 12.090 4.010 ;
        RECT  11.850 1.770 12.090 4.010 ;
        RECT  10.700 3.700 11.140 4.140 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.320 5.600 ;
        RECT  11.770 4.610 12.170 5.600 ;
        RECT  10.540 4.380 10.780 5.600 ;
        RECT  9.170 4.510 9.410 5.600 ;
        RECT  6.450 4.710 6.850 5.600 ;
        RECT  5.260 4.710 5.660 5.600 ;
        RECT  2.340 4.710 2.740 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.320 0.740 ;
        RECT  10.610 0.000 11.550 0.980 ;
        RECT  8.880 0.000 9.280 0.980 ;
        RECT  5.940 0.000 6.180 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.710 ;
        RECT  1.590 3.470 2.430 3.710 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.230 2.190 3.470 3.730 ;
        RECT  4.510 1.660 4.750 3.720 ;
        RECT  5.480 3.220 6.370 3.460 ;
        RECT  4.510 3.400 5.720 3.720 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.740 ;
        RECT  5.010 1.500 6.420 1.740 ;
        RECT  3.900 1.180 4.210 2.000 ;
        RECT  3.690 1.600 4.210 2.000 ;
        RECT  6.180 1.500 6.420 2.500 ;
        RECT  6.180 2.260 6.730 2.500 ;
        RECT  3.970 1.180 4.210 3.730 ;
        RECT  6.710 1.470 6.950 2.020 ;
        RECT  6.710 1.780 7.210 2.020 ;
        RECT  5.700 2.420 5.940 2.980 ;
        RECT  6.970 1.780 7.210 2.980 ;
        RECT  5.700 2.740 7.400 2.980 ;
        RECT  7.160 2.740 7.400 3.730 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 2.390 4.270 ;
        RECT  2.150 4.220 7.270 4.460 ;
        RECT  7.050 4.320 7.980 4.560 ;
        RECT  8.110 1.770 8.720 2.010 ;
        RECT  8.480 1.770 8.720 2.660 ;
        RECT  8.380 2.420 8.620 4.030 ;
        RECT  8.380 3.790 8.960 4.030 ;
        RECT  7.450 1.290 9.380 1.530 ;
        RECT  7.450 1.290 7.690 2.490 ;
        RECT  7.450 2.250 8.140 2.490 ;
        RECT  9.130 1.290 9.380 2.740 ;
        RECT  9.130 2.500 10.380 2.740 ;
        RECT  7.900 2.250 8.140 4.000 ;
        RECT  9.910 1.690 10.900 1.930 ;
        RECT  8.860 3.050 10.900 3.290 ;
        RECT  10.660 1.690 10.900 3.300 ;
        RECT  9.980 3.050 10.900 3.300 ;
        RECT  9.980 3.050 10.220 3.900 ;
    END
END dfcrn2

MACRO dfcrn1
    CLASS CORE ;
    FOREIGN dfcrn1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.020 5.460 2.770 ;
        RECT  5.000 2.500 5.240 3.160 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.031  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.700 3.610 11.610 4.140 ;
        RECT  11.290 1.210 11.530 4.140 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.760 5.600 ;
        RECT  10.720 4.380 10.960 5.600 ;
        RECT  9.420 3.530 9.660 5.600 ;
        RECT  6.450 4.710 6.850 5.600 ;
        RECT  5.260 4.710 5.660 5.600 ;
        RECT  2.350 4.710 2.750 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.760 0.740 ;
        RECT  10.610 0.000 11.010 0.980 ;
        RECT  8.880 0.000 9.280 0.980 ;
        RECT  5.940 0.000 6.180 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.710 ;
        RECT  1.590 3.470 2.430 3.710 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.230 2.190 3.470 3.730 ;
        RECT  4.510 1.660 4.750 3.720 ;
        RECT  5.480 3.220 6.370 3.460 ;
        RECT  4.510 3.400 5.720 3.720 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.740 ;
        RECT  5.010 1.500 6.420 1.740 ;
        RECT  3.900 1.180 4.210 2.000 ;
        RECT  3.690 1.600 4.210 2.000 ;
        RECT  6.180 1.500 6.420 2.500 ;
        RECT  6.180 2.260 6.730 2.500 ;
        RECT  3.970 1.180 4.210 3.730 ;
        RECT  6.710 1.470 6.950 2.020 ;
        RECT  6.710 1.780 7.210 2.020 ;
        RECT  5.700 2.420 5.940 2.980 ;
        RECT  6.970 1.780 7.210 2.980 ;
        RECT  5.700 2.740 7.400 2.980 ;
        RECT  7.160 2.740 7.400 3.730 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 2.390 4.270 ;
        RECT  2.150 4.220 7.270 4.460 ;
        RECT  7.050 4.320 7.980 4.560 ;
        RECT  8.110 1.770 8.720 2.010 ;
        RECT  8.480 1.770 8.720 2.660 ;
        RECT  8.380 2.420 8.620 4.030 ;
        RECT  8.380 3.790 8.960 4.030 ;
        RECT  7.450 1.290 9.380 1.530 ;
        RECT  7.450 1.290 7.690 2.490 ;
        RECT  9.130 1.290 9.380 2.490 ;
        RECT  7.450 2.250 8.140 2.490 ;
        RECT  9.130 2.250 10.540 2.490 ;
        RECT  10.300 2.250 10.540 2.820 ;
        RECT  7.900 2.250 8.140 4.000 ;
        RECT  9.910 1.550 11.050 1.790 ;
        RECT  9.910 1.550 10.310 2.010 ;
        RECT  8.860 3.050 10.220 3.290 ;
        RECT  10.810 1.550 11.050 3.300 ;
        RECT  9.980 3.060 11.050 3.300 ;
        RECT  9.980 3.050 10.220 4.620 ;
    END
END dfcrn1

MACRO dfcrb4
    CLASS CORE ;
    FOREIGN dfcrb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.550 0.980 8.380 1.220 ;
        RECT  5.100 1.510 6.790 1.750 ;
        RECT  6.550 0.980 6.790 1.750 ;
        RECT  5.100 1.460 5.540 1.900 ;
        RECT  5.290 1.460 5.530 2.620 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.340 0.800 2.740 ;
        RECT  0.120 2.340 0.500 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.550 2.740 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.946  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.970 2.020 12.820 2.460 ;
        RECT  12.030 1.070 12.430 2.460 ;
        RECT  11.970 1.420 12.370 3.470 ;
        RECT  10.670 2.700 12.370 3.100 ;
        RECT  10.550 1.420 12.430 1.820 ;
        RECT  10.670 2.700 11.070 3.990 ;
        RECT  10.550 1.070 10.950 1.820 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.867  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.510 1.460 15.390 1.860 ;
        RECT  14.990 1.120 15.390 1.860 ;
        RECT  14.430 2.300 14.830 3.350 ;
        RECT  14.060 1.460 14.500 2.700 ;
        RECT  13.310 2.300 14.830 2.700 ;
        RECT  13.510 1.070 13.910 1.860 ;
        RECT  13.310 2.300 13.710 4.330 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.680 5.600 ;
        RECT  14.060 4.420 14.460 5.600 ;
        RECT  12.740 4.620 13.140 5.600 ;
        RECT  11.410 4.400 11.810 5.600 ;
        RECT  10.070 4.300 10.470 5.600 ;
        RECT  8.810 4.300 9.050 5.600 ;
        RECT  6.040 4.710 6.440 5.600 ;
        RECT  4.620 4.710 5.020 5.600 ;
        RECT  1.990 4.260 2.390 5.600 ;
        RECT  0.720 4.380 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.680 0.740 ;
        RECT  14.250 0.000 14.650 0.980 ;
        RECT  12.770 0.000 13.170 0.980 ;
        RECT  11.290 0.000 11.690 0.980 ;
        RECT  8.620 0.000 9.020 0.890 ;
        RECT  5.690 0.000 6.090 1.260 ;
        RECT  2.030 0.000 2.430 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.850 1.290 2.090 ;
        RECT  1.050 2.520 1.490 2.920 ;
        RECT  1.050 1.850 1.290 3.210 ;
        RECT  0.980 2.970 1.220 3.660 ;
        RECT  0.150 3.420 1.220 3.660 ;
        RECT  2.800 1.680 3.220 2.080 ;
        RECT  2.980 1.680 3.220 3.590 ;
        RECT  2.810 3.350 3.050 3.920 ;
        RECT  1.590 1.140 4.280 1.380 ;
        RECT  1.590 1.140 1.830 2.300 ;
        RECT  1.780 2.060 2.020 3.890 ;
        RECT  1.460 3.650 2.020 3.890 ;
        RECT  4.100 1.740 4.680 1.980 ;
        RECT  4.100 1.740 4.340 3.950 ;
        RECT  4.030 3.550 5.730 3.790 ;
        RECT  4.030 3.550 4.430 3.950 ;
        RECT  3.620 1.680 3.860 3.160 ;
        RECT  6.250 2.840 6.490 3.580 ;
        RECT  5.970 3.340 6.490 3.580 ;
        RECT  3.460 2.920 3.700 4.460 ;
        RECT  5.970 3.340 6.210 4.460 ;
        RECT  3.290 4.220 6.210 4.460 ;
        RECT  3.290 4.220 3.690 4.620 ;
        RECT  5.770 2.000 6.720 2.240 ;
        RECT  6.320 2.000 6.720 2.400 ;
        RECT  6.480 2.360 6.970 2.600 ;
        RECT  4.580 2.220 4.820 3.100 ;
        RECT  5.770 2.000 6.010 3.100 ;
        RECT  4.580 2.860 6.010 3.100 ;
        RECT  6.730 2.360 6.970 4.090 ;
        RECT  7.880 1.940 8.120 3.360 ;
        RECT  7.880 3.120 8.550 3.360 ;
        RECT  8.310 3.120 8.550 4.620 ;
        RECT  7.990 4.380 8.550 4.620 ;
        RECT  7.390 1.460 9.630 1.700 ;
        RECT  7.060 1.880 7.630 2.120 ;
        RECT  9.390 1.460 9.630 2.940 ;
        RECT  9.390 2.700 9.950 2.940 ;
        RECT  7.390 1.460 7.630 4.040 ;
        RECT  7.390 3.640 7.790 4.040 ;
        RECT  9.930 1.390 10.170 2.300 ;
        RECT  9.930 2.060 11.360 2.300 ;
        RECT  10.190 2.060 11.360 2.460 ;
        RECT  8.360 2.560 9.150 2.800 ;
        RECT  8.910 2.560 9.150 3.680 ;
        RECT  10.190 2.060 10.430 3.680 ;
        RECT  8.910 3.440 10.430 3.680 ;
    END
END dfcrb4

MACRO dfcrb2
    CLASS CORE ;
    FOREIGN dfcrb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.020 5.460 2.770 ;
        RECT  5.000 2.500 5.240 3.160 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.318  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.450 3.330 12.260 3.580 ;
        RECT  11.820 3.140 12.260 3.580 ;
        RECT  11.820 1.620 12.060 3.580 ;
        RECT  11.500 1.620 12.060 1.860 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.189  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.880 3.140 13.880 3.650 ;
        RECT  13.490 1.850 13.880 3.650 ;
        RECT  12.880 1.850 13.880 2.090 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 14.000 5.600 ;
        RECT  13.530 4.280 13.770 5.600 ;
        RECT  12.220 4.290 12.460 5.600 ;
        RECT  10.660 4.710 11.060 5.600 ;
        RECT  9.340 4.510 9.580 5.600 ;
        RECT  6.450 4.710 6.850 5.600 ;
        RECT  5.260 4.710 5.660 5.600 ;
        RECT  2.340 4.710 2.740 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 14.000 0.740 ;
        RECT  13.450 0.000 13.850 0.890 ;
        RECT  12.090 0.000 12.490 0.890 ;
        RECT  10.730 0.000 11.130 0.890 ;
        RECT  8.880 0.000 9.280 0.980 ;
        RECT  5.940 0.000 6.180 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.710 ;
        RECT  1.590 3.470 2.430 3.710 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.230 2.190 3.470 3.730 ;
        RECT  4.510 1.660 4.750 3.720 ;
        RECT  5.480 3.220 6.370 3.460 ;
        RECT  4.510 3.400 5.720 3.720 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.740 ;
        RECT  5.010 1.500 6.420 1.740 ;
        RECT  3.900 1.180 4.210 2.000 ;
        RECT  3.690 1.600 4.210 2.000 ;
        RECT  6.180 1.500 6.420 2.500 ;
        RECT  6.180 2.260 6.730 2.500 ;
        RECT  3.970 1.180 4.210 3.730 ;
        RECT  6.710 1.470 6.950 2.020 ;
        RECT  6.710 1.780 7.210 2.020 ;
        RECT  5.700 2.420 5.940 2.980 ;
        RECT  6.970 1.780 7.210 2.980 ;
        RECT  5.700 2.740 7.400 2.980 ;
        RECT  7.160 2.740 7.400 3.730 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 2.390 4.270 ;
        RECT  2.150 4.220 7.300 4.460 ;
        RECT  7.070 4.370 7.980 4.610 ;
        RECT  8.110 1.770 8.720 2.010 ;
        RECT  8.480 1.770 8.720 2.660 ;
        RECT  8.380 2.420 8.620 4.030 ;
        RECT  8.380 3.790 8.960 4.030 ;
        RECT  10.080 1.690 11.080 1.930 ;
        RECT  10.840 2.590 11.550 2.830 ;
        RECT  8.860 3.050 9.760 3.300 ;
        RECT  9.520 3.050 9.760 3.820 ;
        RECT  10.840 1.690 11.080 3.820 ;
        RECT  9.520 3.580 11.080 3.820 ;
        RECT  9.540 1.130 12.620 1.370 ;
        RECT  7.450 1.290 9.780 1.530 ;
        RECT  7.450 1.290 7.690 2.490 ;
        RECT  12.380 1.130 12.620 2.710 ;
        RECT  7.450 2.250 8.140 2.490 ;
        RECT  9.130 1.290 9.380 2.740 ;
        RECT  12.380 2.470 13.030 2.710 ;
        RECT  9.130 2.500 10.450 2.740 ;
        RECT  7.900 2.250 8.140 4.000 ;
    END
END dfcrb2

MACRO dfcrb1
    CLASS CORE ;
    FOREIGN dfcrb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.020 5.460 2.770 ;
        RECT  5.000 2.500 5.240 3.160 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.240  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.020 3.130 11.780 3.370 ;
        RECT  11.540 1.170 11.780 3.370 ;
        RECT  11.260 1.170 11.780 1.900 ;
        RECT  10.950 1.170 11.780 1.410 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.003  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.330 1.540 12.760 3.580 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.880 5.600 ;
        RECT  11.840 4.030 12.080 5.600 ;
        RECT  10.660 4.710 11.060 5.600 ;
        RECT  9.170 4.510 9.410 5.600 ;
        RECT  6.450 4.710 6.850 5.600 ;
        RECT  5.260 4.710 5.660 5.600 ;
        RECT  2.340 4.710 2.740 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.880 0.740 ;
        RECT  11.730 0.000 12.130 0.890 ;
        RECT  8.880 0.000 9.280 0.980 ;
        RECT  5.940 0.000 6.180 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.710 ;
        RECT  1.590 3.470 2.430 3.710 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.230 2.190 3.470 3.730 ;
        RECT  4.510 1.660 4.750 3.720 ;
        RECT  5.480 3.220 6.370 3.460 ;
        RECT  4.510 3.400 5.720 3.720 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.740 ;
        RECT  5.010 1.500 6.420 1.740 ;
        RECT  3.900 1.180 4.210 2.000 ;
        RECT  3.690 1.600 4.210 2.000 ;
        RECT  6.180 1.500 6.420 2.500 ;
        RECT  6.180 2.260 6.730 2.500 ;
        RECT  3.970 1.180 4.210 3.730 ;
        RECT  6.710 1.470 6.950 2.020 ;
        RECT  6.710 1.780 7.210 2.020 ;
        RECT  5.700 2.420 5.940 2.980 ;
        RECT  6.970 1.780 7.210 2.980 ;
        RECT  5.700 2.740 7.400 2.980 ;
        RECT  7.160 2.740 7.400 3.730 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 2.390 4.270 ;
        RECT  2.150 4.220 7.300 4.460 ;
        RECT  7.070 4.370 7.980 4.610 ;
        RECT  8.110 1.770 8.720 2.010 ;
        RECT  8.480 1.770 8.720 2.660 ;
        RECT  8.380 2.420 8.620 4.030 ;
        RECT  8.380 3.790 8.960 4.030 ;
        RECT  7.450 1.290 9.380 1.530 ;
        RECT  7.450 1.290 7.690 2.490 ;
        RECT  9.130 1.290 9.380 2.490 ;
        RECT  7.450 2.250 8.140 2.490 ;
        RECT  9.130 2.250 10.300 2.490 ;
        RECT  10.060 2.250 10.300 2.820 ;
        RECT  7.900 2.250 8.140 4.000 ;
        RECT  9.910 1.690 10.780 1.930 ;
        RECT  10.540 2.590 11.300 2.830 ;
        RECT  8.860 3.050 9.760 3.300 ;
        RECT  9.520 3.050 9.760 3.820 ;
        RECT  10.540 1.690 10.780 3.820 ;
        RECT  9.520 3.580 10.780 3.820 ;
    END
END dfcrb1

MACRO dfcfq4
    CLASS CORE ;
    FOREIGN dfcfq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.580 2.860 10.020 3.580 ;
        RECT  9.400 2.860 10.020 3.260 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.310 2.000 0.560 2.920 ;
        RECT  0.120 2.000 0.560 2.460 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.280 2.020 2.740 2.460 ;
        RECT  2.330 2.020 2.570 3.220 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.632  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.360 1.630 12.820 2.460 ;
        RECT  12.370 1.630 12.770 3.870 ;
        RECT  11.060 3.550 12.770 3.790 ;
        RECT  11.400 1.630 12.820 1.870 ;
        RECT  11.060 3.090 11.300 3.790 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 13.440 5.600 ;
        RECT  12.840 4.620 13.240 5.600 ;
        RECT  11.540 4.620 11.940 5.600 ;
        RECT  10.200 4.620 10.600 5.600 ;
        RECT  8.900 4.620 9.300 5.600 ;
        RECT  5.950 4.710 6.350 5.600 ;
        RECT  4.660 4.620 5.060 5.600 ;
        RECT  1.990 4.380 2.390 5.600 ;
        RECT  0.720 4.440 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 13.440 0.740 ;
        RECT  12.180 0.000 12.580 0.980 ;
        RECT  10.830 0.000 11.230 0.980 ;
        RECT  8.670 0.000 9.070 0.890 ;
        RECT  5.540 0.000 5.940 0.890 ;
        RECT  2.310 0.000 2.710 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.510 1.610 2.040 2.010 ;
        RECT  1.800 1.610 2.040 2.690 ;
        RECT  1.740 2.450 1.980 3.920 ;
        RECT  1.460 3.520 1.980 3.920 ;
        RECT  3.000 1.610 3.240 2.460 ;
        RECT  2.980 2.220 3.220 2.940 ;
        RECT  2.810 2.700 3.050 4.500 ;
        RECT  4.480 1.620 4.720 2.440 ;
        RECT  4.070 2.200 4.720 2.440 ;
        RECT  4.070 2.200 4.310 3.750 ;
        RECT  4.070 3.320 5.740 3.560 ;
        RECT  4.070 3.320 4.470 3.750 ;
        RECT  5.500 3.320 5.740 3.880 ;
        RECT  3.590 1.560 4.060 1.960 ;
        RECT  5.790 2.660 6.230 3.060 ;
        RECT  3.590 1.560 3.830 3.370 ;
        RECT  3.370 3.130 3.610 4.360 ;
        RECT  4.380 4.100 5.400 4.340 ;
        RECT  3.370 4.120 4.620 4.360 ;
        RECT  5.990 2.660 6.230 4.390 ;
        RECT  5.230 4.150 6.230 4.390 ;
        RECT  5.980 1.690 6.620 1.930 ;
        RECT  5.980 1.690 6.220 2.410 ;
        RECT  5.240 2.170 6.710 2.410 ;
        RECT  5.240 2.170 5.480 2.920 ;
        RECT  4.560 2.680 5.480 2.920 ;
        RECT  6.470 2.170 6.710 3.710 ;
        RECT  6.470 3.470 7.040 3.710 ;
        RECT  6.800 3.470 7.040 4.200 ;
        RECT  2.950 0.980 5.310 1.220 ;
        RECT  6.190 0.990 7.190 1.230 ;
        RECT  0.800 1.130 3.190 1.370 ;
        RECT  5.070 1.130 6.430 1.370 ;
        RECT  0.150 1.520 1.040 1.760 ;
        RECT  6.950 0.990 7.190 3.230 ;
        RECT  0.800 2.930 1.500 3.170 ;
        RECT  6.950 2.990 7.520 3.230 ;
        RECT  0.800 1.130 1.040 3.400 ;
        RECT  0.230 3.160 1.040 3.400 ;
        RECT  0.230 3.160 0.470 3.880 ;
        RECT  7.280 2.990 7.520 4.620 ;
        RECT  7.280 4.380 8.220 4.620 ;
        RECT  8.090 1.610 8.490 2.010 ;
        RECT  8.240 1.610 8.480 3.620 ;
        RECT  8.380 3.380 8.620 4.140 ;
        RECT  7.430 1.130 9.680 1.370 ;
        RECT  9.440 1.130 9.680 2.110 ;
        RECT  9.440 1.870 10.260 2.110 ;
        RECT  9.860 1.870 10.260 2.360 ;
        RECT  7.430 1.130 7.670 2.750 ;
        RECT  7.430 2.510 8.000 2.750 ;
        RECT  7.760 2.510 8.000 3.520 ;
        RECT  10.130 1.230 10.820 1.470 ;
        RECT  8.720 2.290 9.120 2.690 ;
        RECT  10.580 2.450 12.070 2.850 ;
        RECT  8.860 2.290 9.100 4.060 ;
        RECT  10.580 1.230 10.820 4.060 ;
        RECT  8.860 3.820 10.820 4.060 ;
    END
END dfcfq4

MACRO dfcfq2
    CLASS CORE ;
    FOREIGN dfcfq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.020 5.460 2.770 ;
        RECT  5.000 2.500 5.240 3.160 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.791  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.230 1.770 12.170 2.170 ;
        RECT  10.700 3.770 12.090 4.010 ;
        RECT  11.850 1.770 12.090 4.010 ;
        RECT  10.700 3.700 11.140 4.140 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.320 5.600 ;
        RECT  11.770 4.610 12.170 5.600 ;
        RECT  10.540 4.380 10.780 5.600 ;
        RECT  9.170 4.510 9.410 5.600 ;
        RECT  6.450 4.710 6.850 5.600 ;
        RECT  5.260 4.710 5.660 5.600 ;
        RECT  2.320 4.710 2.720 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.320 0.740 ;
        RECT  10.610 0.000 11.550 0.980 ;
        RECT  8.880 0.000 9.280 0.980 ;
        RECT  5.940 0.000 6.180 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 1.690 4.270 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.230 2.190 3.470 3.730 ;
        RECT  4.510 1.660 4.750 3.720 ;
        RECT  5.480 3.220 6.370 3.460 ;
        RECT  4.510 3.400 5.720 3.720 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.740 ;
        RECT  5.010 1.500 6.420 1.740 ;
        RECT  3.900 1.180 4.210 2.000 ;
        RECT  3.690 1.600 4.210 2.000 ;
        RECT  6.180 1.500 6.420 2.500 ;
        RECT  6.180 2.260 6.730 2.500 ;
        RECT  3.970 1.180 4.210 3.730 ;
        RECT  6.710 1.470 6.950 2.020 ;
        RECT  6.710 1.780 7.210 2.020 ;
        RECT  5.700 2.420 5.940 2.980 ;
        RECT  6.970 1.780 7.210 2.980 ;
        RECT  5.700 2.740 7.400 2.980 ;
        RECT  7.160 2.740 7.400 3.730 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.630 ;
        RECT  1.590 3.390 2.390 3.630 ;
        RECT  2.150 3.390 2.390 4.460 ;
        RECT  2.150 4.220 7.300 4.460 ;
        RECT  7.070 4.370 7.980 4.610 ;
        RECT  8.110 1.770 8.720 2.010 ;
        RECT  8.480 1.770 8.720 2.660 ;
        RECT  8.380 2.420 8.620 4.030 ;
        RECT  8.380 3.790 8.960 4.030 ;
        RECT  7.450 1.290 9.380 1.530 ;
        RECT  7.450 1.290 7.690 2.490 ;
        RECT  9.130 1.290 9.380 2.490 ;
        RECT  7.450 2.250 8.140 2.490 ;
        RECT  9.130 2.250 10.300 2.490 ;
        RECT  10.060 2.250 10.300 2.820 ;
        RECT  7.900 2.250 8.140 4.000 ;
        RECT  9.910 1.690 10.780 1.930 ;
        RECT  10.540 1.690 10.780 2.620 ;
        RECT  10.540 2.380 11.050 2.620 ;
        RECT  8.860 3.050 9.920 3.300 ;
        RECT  10.810 2.380 11.050 3.300 ;
        RECT  8.860 3.060 11.050 3.300 ;
        RECT  9.980 3.060 10.220 3.900 ;
    END
END dfcfq2

MACRO dfcfq1
    CLASS CORE ;
    FOREIGN dfcfq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.020 5.460 2.770 ;
        RECT  5.000 2.500 5.240 3.160 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.031  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.700 3.610 11.610 4.140 ;
        RECT  11.290 1.210 11.530 4.140 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.760 5.600 ;
        RECT  10.720 4.380 10.960 5.600 ;
        RECT  9.170 4.510 9.410 5.600 ;
        RECT  6.450 4.710 6.850 5.600 ;
        RECT  5.260 4.710 5.660 5.600 ;
        RECT  2.320 4.710 2.720 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.760 0.740 ;
        RECT  10.610 0.000 11.010 0.980 ;
        RECT  8.880 0.000 9.280 0.980 ;
        RECT  5.940 0.000 6.180 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 1.690 4.270 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.230 2.190 3.470 3.730 ;
        RECT  4.510 1.660 4.750 3.720 ;
        RECT  5.480 3.220 6.370 3.460 ;
        RECT  4.510 3.400 5.720 3.720 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.740 ;
        RECT  5.010 1.500 6.420 1.740 ;
        RECT  3.900 1.180 4.210 2.000 ;
        RECT  3.690 1.600 4.210 2.000 ;
        RECT  6.180 1.500 6.420 2.500 ;
        RECT  6.180 2.260 6.730 2.500 ;
        RECT  3.970 1.180 4.210 3.730 ;
        RECT  6.710 1.470 6.950 2.020 ;
        RECT  6.710 1.780 7.210 2.020 ;
        RECT  5.700 2.420 5.940 2.980 ;
        RECT  6.970 1.780 7.210 2.980 ;
        RECT  5.700 2.740 7.400 2.980 ;
        RECT  7.160 2.740 7.400 3.730 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.630 ;
        RECT  1.590 3.390 2.390 3.630 ;
        RECT  2.150 3.390 2.390 4.460 ;
        RECT  2.150 4.220 7.300 4.460 ;
        RECT  7.070 4.370 7.980 4.610 ;
        RECT  8.110 1.770 8.720 2.010 ;
        RECT  8.480 1.770 8.720 2.660 ;
        RECT  8.380 2.420 8.620 4.030 ;
        RECT  8.380 3.790 8.960 4.030 ;
        RECT  7.450 1.290 9.380 1.530 ;
        RECT  7.450 1.290 7.690 2.490 ;
        RECT  9.130 1.290 9.380 2.490 ;
        RECT  7.450 2.250 8.140 2.490 ;
        RECT  9.130 2.250 10.390 2.490 ;
        RECT  10.150 2.250 10.390 2.820 ;
        RECT  7.900 2.250 8.140 4.000 ;
        RECT  10.240 1.550 11.050 1.790 ;
        RECT  9.910 1.690 10.490 1.930 ;
        RECT  8.860 3.050 9.760 3.300 ;
        RECT  10.810 1.550 11.050 3.300 ;
        RECT  10.220 3.060 11.050 3.300 ;
        RECT  9.520 3.050 9.760 3.820 ;
        RECT  10.220 3.060 10.460 3.820 ;
        RECT  9.520 3.580 10.460 3.820 ;
    END
END dfcfq1

MACRO dfcfb4
    CLASS CORE ;
    FOREIGN dfcfb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.560 2.490 6.100 3.020 ;
        RECT  5.300 2.490 6.100 2.890 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.810 3.020 ;
        RECT  0.120 2.490 0.500 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.210 2.020 2.740 2.550 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.716  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 2.970 11.270 3.370 ;
        RECT  9.020 1.530 10.840 1.770 ;
        RECT  9.020 1.530 9.480 3.370 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.718  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.170 2.970 13.880 3.370 ;
        RECT  11.990 1.610 13.750 1.850 ;
        RECT  12.380 1.610 12.820 3.370 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  15.560 4.400 15.960 5.600 ;
        RECT  14.220 4.400 14.620 5.600 ;
        RECT  12.920 4.400 13.320 5.600 ;
        RECT  11.610 4.400 12.010 5.600 ;
        RECT  10.310 4.400 10.710 5.600 ;
        RECT  8.960 4.400 9.360 5.600 ;
        RECT  6.170 4.710 6.570 5.600 ;
        RECT  4.950 4.710 5.350 5.600 ;
        RECT  1.990 4.710 2.390 5.600 ;
        RECT  0.720 4.260 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  13.940 0.000 14.340 0.890 ;
        RECT  12.670 0.000 13.070 0.890 ;
        RECT  11.100 0.000 11.500 0.890 ;
        RECT  9.770 0.000 10.170 0.890 ;
        RECT  8.420 0.000 8.820 0.890 ;
        RECT  5.500 0.000 5.900 1.640 ;
        RECT  1.700 0.000 2.100 0.890 ;
        RECT  0.750 0.000 1.150 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.770 0.550 2.250 ;
        RECT  0.150 2.010 1.080 2.250 ;
        RECT  0.840 2.080 1.410 2.320 ;
        RECT  1.090 2.620 1.490 3.020 ;
        RECT  1.170 2.080 1.410 3.500 ;
        RECT  0.150 3.260 1.410 3.500 ;
        RECT  2.820 1.460 3.220 1.780 ;
        RECT  2.980 1.460 3.220 3.450 ;
        RECT  2.750 3.050 3.220 3.450 ;
        RECT  4.200 1.420 4.700 1.820 ;
        RECT  4.200 1.420 4.440 2.290 ;
        RECT  4.090 2.080 4.330 3.500 ;
        RECT  4.090 3.260 5.990 3.500 ;
        RECT  3.460 1.470 3.960 1.870 ;
        RECT  3.460 1.470 3.700 2.400 ;
        RECT  3.570 2.160 3.810 3.980 ;
        RECT  6.340 2.500 6.580 3.980 ;
        RECT  3.570 3.740 6.580 3.980 ;
        RECT  6.320 1.350 6.560 2.250 ;
        RECT  4.850 2.010 7.060 2.250 ;
        RECT  6.320 2.000 7.060 2.250 ;
        RECT  4.730 2.170 5.080 2.390 ;
        RECT  4.730 2.170 4.970 2.900 ;
        RECT  4.570 2.500 4.970 2.900 ;
        RECT  6.820 2.000 7.060 3.430 ;
        RECT  6.950 3.190 7.190 3.810 ;
        RECT  2.330 0.980 3.730 1.220 ;
        RECT  1.520 1.140 2.570 1.380 ;
        RECT  1.520 1.140 1.970 1.630 ;
        RECT  1.730 1.140 1.970 4.140 ;
        RECT  1.460 3.740 1.970 4.140 ;
        RECT  1.460 3.900 3.020 4.140 ;
        RECT  2.780 3.900 3.020 4.620 ;
        RECT  4.470 4.230 7.330 4.470 ;
        RECT  7.090 4.360 7.780 4.600 ;
        RECT  2.780 4.380 4.720 4.620 ;
        RECT  7.800 1.460 8.040 2.390 ;
        RECT  7.800 2.150 8.530 2.390 ;
        RECT  8.290 2.150 8.530 3.430 ;
        RECT  6.980 1.440 7.540 1.680 ;
        RECT  13.190 2.150 14.130 2.550 ;
        RECT  13.190 2.310 15.470 2.550 ;
        RECT  15.070 2.280 15.470 2.680 ;
        RECT  7.300 1.440 7.540 2.950 ;
        RECT  7.430 2.710 7.670 4.000 ;
        RECT  14.270 2.310 14.510 4.000 ;
        RECT  7.430 3.760 14.510 4.000 ;
        RECT  11.190 1.130 15.570 1.370 ;
        RECT  15.170 1.130 15.570 1.920 ;
        RECT  15.170 1.600 15.950 1.920 ;
        RECT  11.190 1.130 11.430 2.460 ;
        RECT  9.980 2.060 11.460 2.460 ;
        RECT  15.710 1.600 15.950 3.570 ;
        RECT  14.820 3.330 15.950 3.570 ;
    END
END dfcfb4

MACRO dfcfb2
    CLASS CORE ;
    FOREIGN dfcfb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.020 5.460 2.770 ;
        RECT  5.000 2.500 5.240 3.160 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.318  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.450 3.330 12.260 3.580 ;
        RECT  11.820 3.140 12.260 3.580 ;
        RECT  11.820 1.620 12.060 3.580 ;
        RECT  11.500 1.620 12.060 1.860 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.189  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.880 3.140 13.880 3.650 ;
        RECT  13.490 1.850 13.880 3.650 ;
        RECT  12.880 1.850 13.880 2.090 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 14.000 5.600 ;
        RECT  13.530 4.280 13.770 5.600 ;
        RECT  12.220 4.290 12.460 5.600 ;
        RECT  10.660 4.710 11.060 5.600 ;
        RECT  9.340 4.510 9.580 5.600 ;
        RECT  6.450 4.710 6.850 5.600 ;
        RECT  5.260 4.710 5.660 5.600 ;
        RECT  2.560 4.710 2.960 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 14.000 0.740 ;
        RECT  13.450 0.000 13.850 0.890 ;
        RECT  12.090 0.000 12.490 0.890 ;
        RECT  10.730 0.000 11.130 0.890 ;
        RECT  8.880 0.000 9.280 0.980 ;
        RECT  5.940 0.000 6.180 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 1.690 4.270 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.230 2.190 3.470 3.730 ;
        RECT  4.510 1.660 4.750 3.720 ;
        RECT  5.480 3.220 6.370 3.460 ;
        RECT  4.510 3.400 5.720 3.720 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.740 ;
        RECT  5.010 1.500 6.420 1.740 ;
        RECT  3.900 1.180 4.210 2.000 ;
        RECT  3.690 1.600 4.210 2.000 ;
        RECT  6.180 1.500 6.420 2.500 ;
        RECT  6.180 2.260 6.730 2.500 ;
        RECT  3.970 1.180 4.210 3.730 ;
        RECT  6.710 1.470 6.950 2.020 ;
        RECT  6.710 1.780 7.210 2.020 ;
        RECT  5.700 2.420 5.940 2.980 ;
        RECT  6.970 1.780 7.210 2.980 ;
        RECT  5.700 2.740 7.400 2.980 ;
        RECT  7.160 2.740 7.400 3.730 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.630 ;
        RECT  1.590 3.390 2.390 3.630 ;
        RECT  2.150 3.390 2.390 4.460 ;
        RECT  2.150 4.220 7.300 4.460 ;
        RECT  7.070 4.370 7.980 4.610 ;
        RECT  8.110 1.770 8.720 2.010 ;
        RECT  8.480 1.770 8.720 2.660 ;
        RECT  8.380 2.420 8.620 4.030 ;
        RECT  8.380 3.790 8.960 4.030 ;
        RECT  10.080 1.690 11.080 1.930 ;
        RECT  10.840 2.590 11.550 2.830 ;
        RECT  8.860 3.050 9.760 3.300 ;
        RECT  9.520 3.050 9.760 3.820 ;
        RECT  10.840 1.690 11.080 3.820 ;
        RECT  9.520 3.580 11.080 3.820 ;
        RECT  9.540 1.130 12.620 1.370 ;
        RECT  7.450 1.290 9.780 1.530 ;
        RECT  7.450 1.290 7.690 2.490 ;
        RECT  12.380 1.130 12.620 2.710 ;
        RECT  7.450 2.250 8.140 2.490 ;
        RECT  9.130 1.290 9.380 2.740 ;
        RECT  12.380 2.470 13.030 2.710 ;
        RECT  9.130 2.500 10.450 2.740 ;
        RECT  7.900 2.250 8.140 4.000 ;
    END
END dfcfb2

MACRO dfcfb1
    CLASS CORE ;
    FOREIGN dfcfb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.020 5.460 2.770 ;
        RECT  5.000 2.500 5.240 3.160 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.216  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.430 0.790 2.830 ;
        RECT  0.120 2.020 0.500 2.830 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.840 3.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.020 3.130 11.780 3.370 ;
        RECT  11.540 1.170 11.780 3.370 ;
        RECT  11.260 1.170 11.780 1.900 ;
        RECT  10.950 1.170 11.780 1.410 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.003  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.330 1.540 12.760 3.580 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 12.880 5.600 ;
        RECT  11.840 4.030 12.080 5.600 ;
        RECT  10.660 4.710 11.060 5.600 ;
        RECT  9.170 4.510 9.410 5.600 ;
        RECT  6.450 4.710 6.850 5.600 ;
        RECT  5.260 4.710 5.660 5.600 ;
        RECT  2.560 4.710 2.960 5.600 ;
        RECT  0.550 4.050 0.790 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 12.880 0.740 ;
        RECT  11.730 0.000 12.130 0.890 ;
        RECT  8.880 0.000 9.280 0.980 ;
        RECT  5.940 0.000 6.180 1.260 ;
        RECT  2.210 1.660 2.680 2.060 ;
        RECT  2.440 0.000 2.680 2.060 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.270 1.750 ;
        RECT  0.150 3.130 1.270 3.370 ;
        RECT  1.030 1.510 1.270 4.270 ;
        RECT  1.030 4.030 1.690 4.270 ;
        RECT  3.030 1.660 3.270 2.430 ;
        RECT  3.230 2.190 3.470 3.730 ;
        RECT  4.510 1.660 4.750 3.720 ;
        RECT  5.480 3.220 6.370 3.460 ;
        RECT  4.510 3.400 5.720 3.720 ;
        RECT  3.900 1.180 5.250 1.420 ;
        RECT  5.010 1.180 5.250 1.740 ;
        RECT  5.010 1.500 6.420 1.740 ;
        RECT  3.900 1.180 4.210 2.000 ;
        RECT  3.690 1.600 4.210 2.000 ;
        RECT  6.180 1.500 6.420 2.500 ;
        RECT  6.180 2.260 6.730 2.500 ;
        RECT  3.970 1.180 4.210 3.730 ;
        RECT  6.710 1.470 6.950 2.020 ;
        RECT  6.710 1.780 7.210 2.020 ;
        RECT  5.700 2.420 5.940 2.980 ;
        RECT  6.970 1.780 7.210 2.980 ;
        RECT  5.700 2.740 7.400 2.980 ;
        RECT  7.160 2.740 7.400 3.730 ;
        RECT  1.590 0.980 2.140 1.220 ;
        RECT  1.590 0.980 1.830 3.630 ;
        RECT  1.590 3.390 2.390 3.630 ;
        RECT  2.150 3.390 2.390 4.460 ;
        RECT  2.150 4.220 7.300 4.460 ;
        RECT  7.070 4.370 7.980 4.610 ;
        RECT  8.110 1.770 8.720 2.010 ;
        RECT  8.480 1.770 8.720 2.660 ;
        RECT  8.380 2.420 8.620 4.030 ;
        RECT  8.380 3.790 8.960 4.030 ;
        RECT  7.450 1.290 9.380 1.530 ;
        RECT  7.450 1.290 7.690 2.490 ;
        RECT  9.130 1.290 9.380 2.490 ;
        RECT  7.450 2.250 8.140 2.490 ;
        RECT  9.130 2.250 10.300 2.490 ;
        RECT  10.060 2.250 10.300 2.820 ;
        RECT  7.900 2.250 8.140 4.000 ;
        RECT  9.910 1.690 10.780 1.930 ;
        RECT  10.540 2.590 11.300 2.830 ;
        RECT  8.860 3.050 9.760 3.300 ;
        RECT  9.520 3.050 9.760 3.820 ;
        RECT  10.540 1.690 10.780 3.820 ;
        RECT  9.520 3.580 10.780 3.820 ;
    END
END dfcfb1

MACRO dfbrb4
    CLASS CORE ;
    FOREIGN dfbrb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.412  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.580 5.620 3.090 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.270 0.670 2.670 ;
        RECT  0.120 2.270 0.500 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.190 2.580 2.760 3.130 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.868  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.370 1.500 15.250 1.740 ;
        RECT  14.850 1.160 15.250 1.740 ;
        RECT  13.110 3.200 15.200 3.600 ;
        RECT  14.610 1.500 15.200 3.600 ;
        RECT  13.370 1.160 13.770 1.740 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.125  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.330 1.750 18.210 2.120 ;
        RECT  17.810 1.140 18.210 2.120 ;
        RECT  15.770 3.290 17.510 3.690 ;
        RECT  16.860 1.750 17.300 3.690 ;
        RECT  16.330 1.120 16.730 2.120 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.700 2.580 11.140 3.020 ;
        RECT  10.360 2.660 10.780 3.080 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 18.480 5.600 ;
        RECT  17.850 4.240 18.250 5.600 ;
        RECT  16.530 4.240 16.930 5.600 ;
        RECT  15.210 4.240 15.610 5.600 ;
        RECT  13.910 4.240 14.310 5.600 ;
        RECT  12.630 4.150 12.870 5.600 ;
        RECT  11.100 4.690 11.510 5.600 ;
        RECT  9.760 4.330 10.180 5.600 ;
        RECT  6.880 4.330 7.300 5.600 ;
        RECT  4.900 4.490 5.320 5.600 ;
        RECT  2.100 4.490 2.500 5.600 ;
        RECT  0.760 4.130 1.080 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 18.480 0.740 ;
        RECT  17.070 0.000 17.470 1.130 ;
        RECT  15.590 0.000 15.990 1.260 ;
        RECT  14.110 0.000 14.510 1.260 ;
        RECT  12.630 0.000 13.030 1.260 ;
        RECT  10.580 0.000 11.000 1.180 ;
        RECT  5.620 0.000 6.020 1.760 ;
        RECT  2.020 0.000 2.440 0.900 ;
        RECT  0.420 0.000 0.830 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.260 1.010 1.670 1.450 ;
        RECT  0.150 1.390 1.310 1.630 ;
        RECT  1.070 1.210 1.310 3.500 ;
        RECT  0.140 3.260 1.310 3.500 ;
        RECT  2.780 1.620 3.270 2.030 ;
        RECT  3.030 1.620 3.270 3.780 ;
        RECT  2.800 3.380 3.270 3.780 ;
        RECT  3.100 1.040 4.200 1.280 ;
        RECT  2.090 1.140 3.340 1.380 ;
        RECT  2.090 1.140 2.330 2.320 ;
        RECT  1.590 2.080 2.330 2.320 ;
        RECT  1.590 1.700 1.830 3.660 ;
        RECT  4.110 1.610 4.680 1.850 ;
        RECT  4.110 1.610 4.350 3.760 ;
        RECT  5.030 3.370 5.980 3.610 ;
        RECT  4.110 3.520 5.270 3.760 ;
        RECT  7.300 2.610 7.540 3.220 ;
        RECT  3.620 1.550 3.860 4.240 ;
        RECT  7.170 2.970 7.410 4.090 ;
        RECT  6.000 3.850 7.410 4.090 ;
        RECT  3.620 4.000 6.240 4.240 ;
        RECT  7.210 1.500 7.450 2.370 ;
        RECT  4.590 2.100 7.450 2.340 ;
        RECT  6.370 2.130 8.020 2.370 ;
        RECT  4.590 2.100 4.830 3.020 ;
        RECT  7.780 2.130 8.020 3.830 ;
        RECT  6.370 2.100 6.610 3.570 ;
        RECT  7.660 3.430 8.060 3.830 ;
        RECT  7.710 1.080 8.980 1.320 ;
        RECT  8.740 1.080 8.980 2.990 ;
        RECT  9.220 1.550 9.460 3.100 ;
        RECT  9.220 2.860 9.860 3.100 ;
        RECT  9.620 2.860 9.860 3.590 ;
        RECT  9.140 3.350 10.840 3.590 ;
        RECT  7.930 1.650 8.500 1.890 ;
        RECT  8.260 1.650 8.500 3.290 ;
        RECT  8.300 3.150 8.540 4.200 ;
        RECT  11.900 3.690 12.520 3.930 ;
        RECT  12.280 2.520 12.520 3.930 ;
        RECT  8.300 3.850 12.140 4.090 ;
        RECT  8.300 3.800 8.800 4.200 ;
        RECT  11.800 1.690 12.230 2.220 ;
        RECT  9.710 1.790 12.230 2.030 ;
        RECT  11.800 1.980 14.370 2.220 ;
        RECT  9.710 1.790 9.950 2.620 ;
        RECT  11.800 1.690 12.040 3.450 ;
    END
END dfbrb4

MACRO dfbrb2
    CLASS CORE ;
    FOREIGN dfbrb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.670 2.580 12.260 3.030 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.500 0.810 2.740 ;
        RECT  0.140 2.020 0.500 2.740 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.070 1.970 2.740 2.460 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.310 3.140 13.940 3.620 ;
        RECT  13.670 1.330 13.910 3.620 ;
        RECT  13.280 1.330 13.910 1.570 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.870 3.140 15.620 3.620 ;
        RECT  15.180 1.330 15.420 3.620 ;
        RECT  14.760 1.330 15.420 1.570 ;
        RECT  14.870 3.140 15.110 3.960 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.333  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.000 1.460 7.240 2.650 ;
        RECT  6.780 1.460 7.240 1.900 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  15.610 4.340 15.850 5.600 ;
        RECT  14.130 4.340 14.370 5.600 ;
        RECT  12.640 4.340 12.880 5.600 ;
        RECT  11.330 4.340 11.570 5.600 ;
        RECT  10.000 4.340 10.240 5.600 ;
        RECT  6.900 4.660 7.300 5.600 ;
        RECT  5.060 4.660 5.460 5.600 ;
        RECT  2.030 4.660 2.430 5.600 ;
        RECT  0.630 4.070 0.870 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  15.580 0.000 15.820 1.070 ;
        RECT  14.100 0.000 14.340 1.070 ;
        RECT  12.620 0.000 12.860 1.070 ;
        RECT  10.550 0.000 10.790 1.100 ;
        RECT  6.050 0.000 6.290 1.680 ;
        RECT  2.380 0.000 2.620 1.730 ;
        RECT  0.820 0.000 1.060 1.120 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 1.000 2.140 1.240 ;
        RECT  1.590 2.730 2.900 2.970 ;
        RECT  1.590 1.000 1.830 3.450 ;
        RECT  3.140 1.340 3.380 3.910 ;
        RECT  2.800 3.670 3.380 3.910 ;
        RECT  4.850 3.420 6.000 3.660 ;
        RECT  4.850 1.720 5.090 3.720 ;
        RECT  4.280 3.480 5.090 3.720 ;
        RECT  3.980 1.240 5.570 1.480 ;
        RECT  3.980 1.240 4.380 1.740 ;
        RECT  3.620 1.500 4.380 1.740 ;
        RECT  5.330 1.240 5.570 2.570 ;
        RECT  5.330 2.330 6.620 2.570 ;
        RECT  3.620 1.500 3.860 3.800 ;
        RECT  7.560 1.720 7.960 2.040 ;
        RECT  5.480 2.890 6.740 3.130 ;
        RECT  7.720 1.720 7.960 3.680 ;
        RECT  6.340 2.890 6.740 3.680 ;
        RECT  7.720 3.280 8.110 3.680 ;
        RECT  6.340 3.360 8.110 3.680 ;
        RECT  0.150 1.540 1.350 1.780 ;
        RECT  0.150 3.130 1.350 3.370 ;
        RECT  1.110 1.540 1.350 4.420 ;
        RECT  7.350 4.140 8.470 4.380 ;
        RECT  1.110 4.180 7.670 4.420 ;
        RECT  9.120 1.720 9.360 2.340 ;
        RECT  9.250 2.100 9.490 3.620 ;
        RECT  9.250 3.220 9.710 3.620 ;
        RECT  9.250 3.300 10.950 3.620 ;
        RECT  11.810 1.310 12.660 1.550 ;
        RECT  12.420 1.310 12.660 2.130 ;
        RECT  12.420 1.890 13.430 2.130 ;
        RECT  10.300 2.770 11.430 3.010 ;
        RECT  11.190 2.770 11.430 3.620 ;
        RECT  12.500 1.890 12.740 3.620 ;
        RECT  11.190 3.380 12.740 3.620 ;
        RECT  8.300 1.240 9.970 1.480 ;
        RECT  8.300 1.240 8.760 1.780 ;
        RECT  9.730 1.240 9.970 2.080 ;
        RECT  9.730 1.840 11.960 2.080 ;
        RECT  8.520 1.240 8.760 3.680 ;
        RECT  8.450 3.280 9.010 3.680 ;
        RECT  8.770 3.280 9.010 4.100 ;
        RECT  14.350 2.690 14.590 4.100 ;
        RECT  8.770 3.860 14.590 4.100 ;
    END
END dfbrb2

MACRO dfbrb1
    CLASS CORE ;
    FOREIGN dfbrb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.670 2.580 12.260 3.030 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.500 0.810 2.740 ;
        RECT  0.140 2.020 0.500 2.740 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.070 1.970 2.740 2.460 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.068  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.260 3.130 14.020 3.580 ;
        RECT  13.780 1.860 14.020 3.580 ;
        RECT  13.270 1.860 14.020 2.100 ;
        RECT  13.270 1.080 13.510 2.100 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.003  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.570 1.560 15.000 3.450 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.333  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.000 1.460 7.240 2.650 ;
        RECT  6.780 1.460 7.240 1.900 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.120 5.600 ;
        RECT  14.080 4.030 14.320 5.600 ;
        RECT  12.730 4.580 13.130 5.600 ;
        RECT  11.330 4.340 11.570 5.600 ;
        RECT  10.000 4.340 10.240 5.600 ;
        RECT  6.900 4.660 7.300 5.600 ;
        RECT  5.060 4.660 5.460 5.600 ;
        RECT  2.030 4.660 2.430 5.600 ;
        RECT  0.630 4.070 0.870 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.120 0.740 ;
        RECT  13.970 0.000 14.370 0.890 ;
        RECT  10.550 0.000 10.790 1.100 ;
        RECT  6.050 0.000 6.290 1.680 ;
        RECT  2.380 0.000 2.620 1.730 ;
        RECT  0.820 0.000 1.060 1.120 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 1.000 2.140 1.240 ;
        RECT  1.590 2.730 2.900 2.970 ;
        RECT  1.590 1.000 1.830 3.450 ;
        RECT  3.140 1.340 3.380 3.910 ;
        RECT  2.800 3.670 3.380 3.910 ;
        RECT  4.850 3.420 6.000 3.660 ;
        RECT  4.850 1.720 5.090 3.720 ;
        RECT  4.280 3.480 5.090 3.720 ;
        RECT  3.980 1.240 5.570 1.480 ;
        RECT  3.980 1.240 4.380 1.740 ;
        RECT  3.620 1.500 4.380 1.740 ;
        RECT  5.330 1.240 5.570 2.570 ;
        RECT  5.330 2.330 6.620 2.570 ;
        RECT  3.620 1.500 3.860 3.800 ;
        RECT  7.560 1.720 7.960 2.120 ;
        RECT  5.480 2.890 6.740 3.130 ;
        RECT  7.720 1.720 7.960 3.680 ;
        RECT  6.340 2.890 6.740 3.680 ;
        RECT  7.720 3.280 8.110 3.680 ;
        RECT  6.340 3.360 8.110 3.680 ;
        RECT  0.150 1.540 1.350 1.780 ;
        RECT  0.150 3.130 1.350 3.370 ;
        RECT  1.110 1.540 1.350 4.420 ;
        RECT  7.350 4.140 8.470 4.380 ;
        RECT  1.110 4.180 7.670 4.420 ;
        RECT  9.120 1.720 9.360 2.340 ;
        RECT  9.250 2.100 9.490 3.620 ;
        RECT  9.250 3.220 9.710 3.620 ;
        RECT  9.250 3.300 10.950 3.620 ;
        RECT  8.300 1.240 9.970 1.480 ;
        RECT  8.300 1.240 8.770 1.780 ;
        RECT  9.730 1.240 9.970 2.080 ;
        RECT  9.730 1.840 11.960 2.080 ;
        RECT  8.530 1.240 8.770 3.680 ;
        RECT  11.870 1.310 12.950 1.550 ;
        RECT  12.710 2.590 13.540 2.830 ;
        RECT  10.300 2.770 11.430 3.010 ;
        RECT  11.190 2.770 11.430 3.730 ;
        RECT  12.710 1.310 12.950 3.730 ;
        RECT  11.190 3.490 12.950 3.730 ;
    END
END dfbrb1

MACRO dfbfb4
    CLASS CORE ;
    FOREIGN dfbfb4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 2.480 6.190 3.020 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.436  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.300 0.800 2.700 ;
        RECT  0.120 2.300 0.500 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 2.210 2.740 3.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.890  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.840 1.660 18.730 1.900 ;
        RECT  17.980 1.660 18.420 3.050 ;
        RECT  16.540 3.050 18.250 3.450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.937  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.830 1.750 15.710 1.990 ;
        RECT  13.920 3.080 15.640 3.320 ;
        RECT  14.620 1.750 15.060 3.320 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.781  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.690 2.790 11.930 3.990 ;
        RECT  11.510 2.460 11.750 3.030 ;
        RECT  8.980 3.750 11.930 3.990 ;
        RECT  6.550 3.760 9.220 4.000 ;
        RECT  6.550 2.540 7.240 3.020 ;
        RECT  6.550 2.540 6.790 4.000 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.040 5.600 ;
        RECT  18.410 4.620 18.810 5.600 ;
        RECT  17.110 4.450 17.510 5.600 ;
        RECT  15.800 4.450 16.200 5.600 ;
        RECT  14.500 4.460 14.900 5.600 ;
        RECT  13.170 4.040 13.570 5.600 ;
        RECT  11.840 4.710 12.240 5.600 ;
        RECT  10.470 4.710 10.870 5.600 ;
        RECT  7.620 4.320 7.860 5.600 ;
        RECT  6.080 4.320 6.480 5.600 ;
        RECT  4.720 4.570 5.120 5.600 ;
        RECT  2.220 4.710 2.620 5.600 ;
        RECT  0.920 4.710 1.320 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.040 0.740 ;
        RECT  17.590 0.000 17.990 1.420 ;
        RECT  16.080 0.000 16.480 0.890 ;
        RECT  14.570 0.000 14.970 1.490 ;
        RECT  11.730 0.000 12.130 0.890 ;
        RECT  6.160 0.000 6.560 1.280 ;
        RECT  2.170 0.000 2.570 0.890 ;
        RECT  0.740 0.000 1.140 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.820 1.280 2.060 ;
        RECT  1.040 2.410 1.480 2.810 ;
        RECT  1.040 1.820 1.280 3.180 ;
        RECT  0.760 2.940 1.280 3.180 ;
        RECT  0.760 2.940 1.000 3.500 ;
        RECT  0.150 3.260 1.000 3.500 ;
        RECT  2.950 1.370 3.190 1.970 ;
        RECT  2.980 1.730 3.220 2.760 ;
        RECT  3.210 2.520 3.450 3.640 ;
        RECT  2.810 3.400 3.450 3.640 ;
        RECT  1.800 1.110 2.040 1.670 ;
        RECT  1.590 1.430 1.830 2.190 ;
        RECT  1.740 1.950 1.980 3.290 ;
        RECT  1.530 3.050 1.770 4.210 ;
        RECT  1.530 3.970 3.790 4.210 ;
        RECT  3.550 3.970 3.790 4.620 ;
        RECT  3.550 4.380 4.340 4.620 ;
        RECT  4.410 1.470 4.990 1.710 ;
        RECT  4.410 1.470 4.650 3.550 ;
        RECT  4.410 3.310 5.890 3.550 ;
        RECT  4.510 3.310 4.750 4.090 ;
        RECT  4.190 3.850 4.750 4.090 ;
        RECT  3.690 0.980 5.780 1.220 ;
        RECT  7.370 1.140 8.390 1.380 ;
        RECT  5.540 0.980 5.780 1.760 ;
        RECT  7.070 1.280 7.610 1.520 ;
        RECT  5.540 1.520 7.310 1.760 ;
        RECT  3.690 0.980 3.930 3.450 ;
        RECT  7.920 1.680 8.160 2.240 ;
        RECT  4.970 2.000 8.620 2.240 ;
        RECT  7.740 2.480 8.620 2.720 ;
        RECT  4.970 2.000 5.210 2.800 ;
        RECT  7.740 2.480 7.990 3.500 ;
        RECT  7.030 3.260 7.990 3.500 ;
        RECT  8.380 2.000 8.620 3.510 ;
        RECT  9.810 1.490 10.440 1.730 ;
        RECT  10.200 1.490 10.440 3.510 ;
        RECT  9.780 3.190 10.440 3.430 ;
        RECT  10.200 3.270 11.450 3.510 ;
        RECT  12.150 2.150 12.550 2.550 ;
        RECT  9.880 4.230 12.410 4.470 ;
        RECT  12.170 2.150 12.410 4.470 ;
        RECT  8.100 4.380 10.120 4.620 ;
        RECT  9.150 0.980 11.270 1.220 ;
        RECT  12.600 0.980 13.860 1.220 ;
        RECT  11.030 1.180 12.840 1.420 ;
        RECT  9.150 0.980 9.390 2.750 ;
        RECT  9.120 2.450 9.360 3.510 ;
        RECT  11.660 1.670 13.500 1.910 ;
        RECT  13.100 1.620 13.500 2.020 ;
        RECT  11.660 1.670 11.900 2.210 ;
        RECT  11.020 1.970 11.900 2.210 ;
        RECT  11.020 1.970 11.260 2.500 ;
        RECT  10.700 2.260 11.260 2.500 ;
        RECT  15.960 2.270 17.510 2.670 ;
        RECT  13.240 1.620 13.480 3.060 ;
        RECT  12.650 2.820 13.480 3.060 ;
        RECT  12.650 2.820 12.890 3.800 ;
        RECT  12.650 3.560 14.680 3.800 ;
        RECT  14.440 3.560 14.680 4.190 ;
        RECT  15.960 2.270 16.200 4.190 ;
        RECT  14.440 3.950 16.200 4.190 ;
    END
END dfbfb4

MACRO dfbfb2
    CLASS CORE ;
    FOREIGN dfbfb2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.670 2.580 12.260 3.030 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.500 0.810 2.740 ;
        RECT  0.140 2.020 0.500 2.740 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.070 1.970 2.740 2.460 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.310 3.140 13.940 3.620 ;
        RECT  13.670 1.330 13.910 3.620 ;
        RECT  13.280 1.330 13.910 1.570 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.870 3.140 15.620 3.620 ;
        RECT  15.180 1.330 15.420 3.620 ;
        RECT  14.760 1.330 15.420 1.570 ;
        RECT  14.870 3.140 15.110 3.960 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.333  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.000 1.460 7.240 2.650 ;
        RECT  6.780 1.460 7.240 1.900 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  15.610 4.340 15.850 5.600 ;
        RECT  14.130 4.340 14.370 5.600 ;
        RECT  12.640 4.340 12.880 5.600 ;
        RECT  11.330 4.340 11.570 5.600 ;
        RECT  10.000 4.340 10.240 5.600 ;
        RECT  6.900 4.660 7.300 5.600 ;
        RECT  5.060 4.660 5.460 5.600 ;
        RECT  2.030 4.660 2.430 5.600 ;
        RECT  0.630 4.070 0.870 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  15.580 0.000 15.820 1.070 ;
        RECT  14.100 0.000 14.340 1.070 ;
        RECT  12.620 0.000 12.860 1.070 ;
        RECT  10.550 0.000 10.790 1.100 ;
        RECT  6.050 0.000 6.290 1.680 ;
        RECT  2.380 0.000 2.620 1.730 ;
        RECT  0.820 0.000 1.060 1.120 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.350 1.780 ;
        RECT  0.150 3.130 1.350 3.370 ;
        RECT  1.110 1.540 1.350 4.420 ;
        RECT  1.110 4.180 1.670 4.420 ;
        RECT  3.140 1.340 3.380 3.910 ;
        RECT  2.800 3.670 3.380 3.910 ;
        RECT  4.850 3.420 6.000 3.660 ;
        RECT  4.850 1.720 5.090 3.720 ;
        RECT  4.280 3.480 5.090 3.720 ;
        RECT  3.980 1.240 5.570 1.480 ;
        RECT  3.980 1.240 4.380 1.740 ;
        RECT  3.620 1.500 4.380 1.740 ;
        RECT  5.330 1.240 5.570 2.570 ;
        RECT  5.330 2.330 6.620 2.570 ;
        RECT  3.620 1.500 3.860 3.800 ;
        RECT  7.560 1.720 7.960 2.120 ;
        RECT  5.480 2.890 6.740 3.130 ;
        RECT  7.720 1.720 7.960 3.680 ;
        RECT  6.340 2.890 6.740 3.680 ;
        RECT  7.720 3.280 8.110 3.680 ;
        RECT  6.340 3.360 8.110 3.680 ;
        RECT  1.590 1.000 2.140 1.240 ;
        RECT  1.590 1.000 1.830 3.860 ;
        RECT  1.590 3.620 2.320 3.860 ;
        RECT  2.080 3.620 2.320 4.420 ;
        RECT  7.350 4.140 8.470 4.380 ;
        RECT  2.080 4.180 7.670 4.420 ;
        RECT  9.120 1.720 9.360 2.340 ;
        RECT  9.250 2.100 9.490 3.620 ;
        RECT  9.250 3.220 9.710 3.620 ;
        RECT  9.250 3.300 10.950 3.620 ;
        RECT  11.810 1.310 12.660 1.550 ;
        RECT  12.420 1.310 12.660 2.130 ;
        RECT  12.420 1.890 13.430 2.130 ;
        RECT  10.300 2.770 11.430 3.010 ;
        RECT  11.190 2.770 11.430 3.620 ;
        RECT  12.500 1.890 12.740 3.620 ;
        RECT  11.190 3.380 12.740 3.620 ;
        RECT  8.300 1.240 9.970 1.480 ;
        RECT  8.300 1.240 8.770 1.780 ;
        RECT  9.730 1.240 9.970 2.080 ;
        RECT  9.730 1.840 11.960 2.080 ;
        RECT  8.530 3.660 9.010 3.900 ;
        RECT  8.530 1.240 8.770 3.900 ;
        RECT  14.350 2.690 14.590 4.100 ;
        RECT  8.710 3.860 14.590 4.100 ;
    END
END dfbfb2

MACRO dfbfb1
    CLASS CORE ;
    FOREIGN dfbfb1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.670 2.580 12.260 3.030 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.500 0.810 2.740 ;
        RECT  0.140 2.020 0.500 2.740 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.070 1.970 2.740 2.460 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.068  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.260 3.130 14.020 3.580 ;
        RECT  13.780 1.860 14.020 3.580 ;
        RECT  13.270 1.860 14.020 2.100 ;
        RECT  13.270 1.080 13.510 2.100 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.003  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.570 1.560 15.000 3.450 ;
        END
    END QN
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.333  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.000 1.460 7.240 2.650 ;
        RECT  6.780 1.460 7.240 1.900 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.120 5.600 ;
        RECT  14.080 4.030 14.320 5.600 ;
        RECT  12.730 4.580 13.130 5.600 ;
        RECT  11.330 4.340 11.570 5.600 ;
        RECT  10.000 4.340 10.240 5.600 ;
        RECT  6.900 4.660 7.300 5.600 ;
        RECT  5.060 4.660 5.460 5.600 ;
        RECT  2.030 4.660 2.430 5.600 ;
        RECT  0.630 4.070 0.870 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.120 0.740 ;
        RECT  13.970 0.000 14.370 0.890 ;
        RECT  10.550 0.000 10.790 1.100 ;
        RECT  6.050 0.000 6.290 1.680 ;
        RECT  2.380 0.000 2.620 1.730 ;
        RECT  0.820 0.000 1.060 1.120 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.350 1.780 ;
        RECT  0.150 3.130 1.350 3.370 ;
        RECT  1.110 1.540 1.350 4.420 ;
        RECT  1.110 4.180 1.670 4.420 ;
        RECT  3.140 1.340 3.380 3.910 ;
        RECT  2.800 3.670 3.380 3.910 ;
        RECT  4.850 3.420 6.000 3.660 ;
        RECT  4.850 1.720 5.090 3.720 ;
        RECT  4.280 3.480 5.090 3.720 ;
        RECT  3.980 1.240 5.570 1.480 ;
        RECT  3.980 1.240 4.380 1.740 ;
        RECT  3.620 1.500 4.380 1.740 ;
        RECT  5.330 1.240 5.570 2.570 ;
        RECT  5.330 2.330 6.620 2.570 ;
        RECT  3.620 1.500 3.860 3.800 ;
        RECT  7.560 1.720 7.960 2.120 ;
        RECT  5.480 2.890 6.740 3.130 ;
        RECT  7.720 1.720 7.960 3.680 ;
        RECT  6.340 2.890 6.740 3.680 ;
        RECT  7.720 3.280 8.110 3.680 ;
        RECT  6.340 3.360 8.110 3.680 ;
        RECT  1.590 1.000 2.140 1.240 ;
        RECT  1.590 1.000 1.830 3.860 ;
        RECT  1.590 3.620 2.320 3.860 ;
        RECT  2.080 3.620 2.320 4.420 ;
        RECT  7.350 4.140 8.470 4.380 ;
        RECT  2.080 4.180 7.670 4.420 ;
        RECT  9.120 1.720 9.360 2.340 ;
        RECT  9.250 2.100 9.490 3.620 ;
        RECT  9.250 3.220 9.710 3.620 ;
        RECT  9.250 3.300 10.950 3.620 ;
        RECT  8.300 1.240 9.970 1.480 ;
        RECT  8.300 1.240 8.770 1.780 ;
        RECT  9.730 1.240 9.970 2.080 ;
        RECT  9.730 1.840 11.960 2.080 ;
        RECT  8.530 1.240 8.770 3.680 ;
        RECT  11.870 1.310 12.950 1.550 ;
        RECT  12.710 2.590 13.540 2.830 ;
        RECT  10.300 2.770 11.430 3.010 ;
        RECT  11.190 2.770 11.430 3.730 ;
        RECT  12.710 1.310 12.950 3.730 ;
        RECT  11.190 3.490 12.950 3.730 ;
    END
END dfbfb1

MACRO deprq4
    CLASS CORE ;
    FOREIGN deprq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.700 2.020 11.190 2.520 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.393  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.740 3.020 ;
        RECT  2.230 2.330 2.630 2.730 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.320 0.780 2.720 ;
        RECT  0.120 2.320 0.500 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.860  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.900 2.920 10.270 3.160 ;
        RECT  10.030 1.510 10.270 3.160 ;
        RECT  8.400 1.880 10.270 2.120 ;
        RECT  9.800 1.510 10.270 2.120 ;
        RECT  8.400 1.510 8.640 2.120 ;
        RECT  7.900 2.860 8.340 3.300 ;
        END
    END Q
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.451  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.580 5.610 3.110 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.720 5.600 ;
        RECT  19.050 4.270 19.450 5.600 ;
        RECT  10.150 4.400 10.550 5.600 ;
        RECT  8.850 4.400 9.250 5.600 ;
        RECT  7.550 4.400 7.950 5.600 ;
        RECT  6.150 4.380 6.550 5.600 ;
        RECT  4.840 4.400 5.240 5.600 ;
        RECT  2.240 3.490 2.480 5.600 ;
        RECT  0.720 4.110 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.720 0.740 ;
        RECT  18.380 0.000 18.780 0.900 ;
        RECT  12.060 0.000 12.300 1.640 ;
        RECT  10.540 0.000 10.940 1.640 ;
        RECT  9.060 0.000 9.460 1.640 ;
        RECT  7.580 0.000 7.980 1.640 ;
        RECT  4.910 0.000 5.310 0.890 ;
        RECT  1.730 0.000 2.130 0.910 ;
        RECT  0.740 0.000 1.140 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.780 1.260 2.020 ;
        RECT  1.020 2.490 1.480 2.890 ;
        RECT  1.020 1.780 1.260 3.510 ;
        RECT  0.150 3.270 1.260 3.510 ;
        RECT  2.800 1.640 3.220 2.040 ;
        RECT  2.980 1.640 3.220 4.590 ;
        RECT  2.730 4.190 3.220 4.590 ;
        RECT  2.390 1.060 4.190 1.300 ;
        RECT  1.590 1.220 2.630 1.460 ;
        RECT  1.590 1.220 1.830 2.250 ;
        RECT  1.730 2.010 1.970 3.370 ;
        RECT  1.540 3.130 1.780 3.800 ;
        RECT  4.400 1.780 4.640 3.650 ;
        RECT  4.070 3.410 4.640 3.650 ;
        RECT  4.520 1.130 5.320 1.370 ;
        RECT  5.080 1.130 5.320 1.950 ;
        RECT  5.080 1.710 6.540 1.950 ;
        RECT  5.860 1.710 6.100 3.660 ;
        RECT  5.410 3.420 6.100 3.660 ;
        RECT  5.880 1.010 7.160 1.250 ;
        RECT  6.920 2.360 9.510 2.600 ;
        RECT  6.920 1.010 7.160 3.650 ;
        RECT  6.720 3.250 7.160 3.650 ;
        RECT  11.280 1.420 11.810 1.780 ;
        RECT  11.570 1.420 11.810 3.120 ;
        RECT  10.890 2.880 11.810 3.120 ;
        RECT  12.540 1.380 13.120 1.620 ;
        RECT  12.540 1.380 12.780 2.660 ;
        RECT  12.240 2.260 12.780 2.660 ;
        RECT  12.240 2.260 12.480 3.210 ;
        RECT  3.550 1.570 3.980 1.970 ;
        RECT  13.500 1.470 13.740 2.100 ;
        RECT  13.020 1.860 13.740 2.100 ;
        RECT  13.020 1.860 13.260 4.140 ;
        RECT  3.550 3.900 13.260 4.140 ;
        RECT  3.550 1.570 3.790 4.500 ;
        RECT  12.660 3.900 13.060 4.520 ;
        RECT  15.250 0.980 16.660 1.220 ;
        RECT  16.420 0.980 16.660 2.310 ;
        RECT  15.940 2.070 16.660 2.310 ;
        RECT  15.940 2.070 16.180 3.170 ;
        RECT  15.600 2.930 16.180 3.170 ;
        RECT  15.460 1.460 16.000 1.830 ;
        RECT  15.460 1.460 15.700 2.690 ;
        RECT  14.940 2.450 15.700 2.690 ;
        RECT  17.310 2.970 17.620 3.170 ;
        RECT  17.380 2.240 17.620 3.170 ;
        RECT  16.900 3.030 17.530 3.270 ;
        RECT  14.940 2.450 15.180 3.660 ;
        RECT  16.900 3.030 17.140 3.660 ;
        RECT  14.940 3.420 17.140 3.660 ;
        RECT  16.900 0.980 17.720 1.220 ;
        RECT  16.900 1.480 17.480 1.880 ;
        RECT  16.900 0.980 17.140 2.790 ;
        RECT  16.420 2.550 17.140 2.790 ;
        RECT  16.420 2.550 16.660 3.160 ;
        RECT  14.980 1.470 15.220 2.210 ;
        RECT  14.460 1.970 15.220 2.210 ;
        RECT  17.860 1.470 18.100 3.880 ;
        RECT  14.460 1.970 14.700 3.520 ;
        RECT  14.070 3.120 14.700 3.520 ;
        RECT  17.730 3.480 18.130 3.880 ;
        RECT  17.380 3.640 18.130 3.880 ;
        RECT  14.070 3.120 14.390 4.140 ;
        RECT  17.380 3.640 17.620 4.140 ;
        RECT  14.070 3.900 17.620 4.140 ;
        RECT  13.980 1.490 14.560 1.730 ;
        RECT  13.980 1.490 14.220 2.580 ;
        RECT  13.530 2.340 14.220 2.580 ;
        RECT  13.530 2.340 13.770 4.620 ;
        RECT  17.920 4.120 18.320 4.620 ;
        RECT  13.530 4.380 18.320 4.620 ;
        RECT  18.340 2.010 18.580 3.180 ;
        RECT  19.160 1.470 19.400 3.180 ;
        RECT  18.340 2.780 19.400 3.180 ;
        RECT  18.340 2.860 20.360 3.180 ;
        RECT  19.960 2.860 20.360 3.450 ;
    END
END deprq4

MACRO deprq2
    CLASS CORE ;
    FOREIGN deprq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.203  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.100 5.620 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.150 4.380 3.860 4.620 ;
        RECT  3.420 3.700 3.860 4.620 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.170 0.550 2.600 ;
        RECT  0.120 1.460 0.500 2.600 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.152  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.250 3.130 16.740 3.580 ;
        RECT  16.250 1.620 16.490 3.580 ;
        END
    END Q
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.500 2.020 13.970 2.490 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.360 5.600 ;
        RECT  16.870 4.170 17.110 5.600 ;
        RECT  15.560 3.190 15.800 5.600 ;
        RECT  14.290 4.400 14.530 5.600 ;
        RECT  12.810 4.400 13.050 5.600 ;
        RECT  10.610 4.650 11.010 5.600 ;
        RECT  9.250 4.650 9.650 5.600 ;
        RECT  5.570 4.610 5.970 5.600 ;
        RECT  4.460 4.610 4.860 5.600 ;
        RECT  1.670 4.300 1.910 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.360 0.740 ;
        RECT  16.810 0.000 17.210 0.890 ;
        RECT  15.510 0.000 15.750 1.460 ;
        RECT  13.980 0.000 14.220 1.290 ;
        RECT  9.340 0.000 9.580 2.110 ;
        RECT  5.570 0.000 5.970 0.890 ;
        RECT  4.280 0.000 4.680 0.890 ;
        RECT  1.770 0.000 2.170 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 2.570 1.500 2.810 ;
        RECT  0.820 1.610 1.060 3.450 ;
        RECT  2.290 1.530 2.530 3.460 ;
        RECT  0.850 0.980 1.540 1.220 ;
        RECT  1.300 0.980 1.540 1.800 ;
        RECT  1.300 1.560 2.030 1.800 ;
        RECT  1.790 1.560 2.030 4.000 ;
        RECT  0.930 3.760 3.140 4.000 ;
        RECT  0.930 3.760 1.170 4.610 ;
        RECT  3.690 1.610 4.260 1.850 ;
        RECT  4.020 1.610 4.260 3.380 ;
        RECT  3.690 3.140 4.260 3.380 ;
        RECT  4.980 1.620 6.100 1.860 ;
        RECT  5.860 2.170 6.310 2.570 ;
        RECT  5.860 1.620 6.100 3.720 ;
        RECT  4.980 3.480 6.100 3.720 ;
        RECT  6.340 1.610 6.880 1.930 ;
        RECT  6.640 1.610 6.880 3.720 ;
        RECT  6.640 2.710 6.910 3.720 ;
        RECT  6.340 3.480 6.910 3.720 ;
        RECT  3.030 1.130 7.360 1.370 ;
        RECT  7.120 1.130 7.360 2.340 ;
        RECT  7.230 2.100 7.470 3.450 ;
        RECT  3.030 1.130 3.270 3.460 ;
        RECT  8.530 1.770 8.920 2.090 ;
        RECT  8.530 1.770 8.770 3.450 ;
        RECT  8.530 3.130 9.060 3.450 ;
        RECT  7.780 1.770 8.230 2.090 ;
        RECT  7.990 1.770 8.230 3.930 ;
        RECT  10.580 2.520 10.820 3.930 ;
        RECT  7.990 3.690 10.820 3.930 ;
        RECT  10.100 1.850 11.300 2.090 ;
        RECT  9.010 2.380 10.340 2.620 ;
        RECT  11.060 1.850 11.300 3.370 ;
        RECT  11.060 3.130 11.860 3.370 ;
        RECT  10.100 1.850 10.340 3.450 ;
        RECT  12.210 1.850 13.260 2.090 ;
        RECT  13.020 1.850 13.260 4.160 ;
        RECT  4.500 2.520 4.740 4.200 ;
        RECT  11.210 3.920 13.790 4.160 ;
        RECT  4.500 3.960 6.580 4.200 ;
        RECT  11.210 3.920 11.450 4.410 ;
        RECT  6.340 4.170 11.450 4.410 ;
        RECT  13.550 3.920 13.790 4.570 ;
        RECT  11.540 1.370 13.740 1.610 ;
        RECT  13.500 1.540 14.450 1.780 ;
        RECT  14.210 1.540 14.450 2.470 ;
        RECT  14.210 2.230 15.020 2.470 ;
        RECT  11.540 1.370 11.780 2.890 ;
        RECT  11.540 2.650 12.520 2.890 ;
        RECT  12.280 2.650 12.520 3.450 ;
        RECT  14.690 1.700 15.940 1.940 ;
        RECT  14.950 2.710 15.940 2.950 ;
        RECT  15.700 1.700 15.940 2.950 ;
        RECT  13.500 2.850 15.190 3.090 ;
        RECT  14.950 2.710 15.190 4.220 ;
    END
END deprq2

MACRO deprq1
    CLASS CORE ;
    FOREIGN deprq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.203  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.100 5.620 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.094  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.150 4.380 3.860 4.620 ;
        RECT  3.420 3.700 3.860 4.620 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.170 0.550 2.600 ;
        RECT  0.120 1.460 0.500 2.600 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.061  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 3.140 16.640 3.580 ;
        RECT  16.320 1.400 16.640 3.580 ;
        END
    END Q
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.500 2.020 13.990 2.490 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  15.750 4.070 15.990 5.600 ;
        RECT  14.390 4.400 14.630 5.600 ;
        RECT  12.910 4.400 13.150 5.600 ;
        RECT  10.610 4.650 11.010 5.600 ;
        RECT  9.250 4.650 9.650 5.600 ;
        RECT  5.570 4.610 5.970 5.600 ;
        RECT  4.460 4.610 4.860 5.600 ;
        RECT  1.670 4.300 1.910 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  15.580 0.000 15.820 1.240 ;
        RECT  13.980 0.000 14.220 1.290 ;
        RECT  9.340 0.000 9.580 2.110 ;
        RECT  5.570 0.000 5.970 0.890 ;
        RECT  4.280 0.000 4.680 0.890 ;
        RECT  1.770 0.000 2.170 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 2.570 1.500 2.810 ;
        RECT  0.820 1.610 1.060 3.450 ;
        RECT  2.290 1.530 2.530 3.460 ;
        RECT  0.850 0.980 1.540 1.220 ;
        RECT  1.300 0.980 1.540 1.800 ;
        RECT  1.300 1.560 2.030 1.800 ;
        RECT  1.790 1.560 2.030 4.000 ;
        RECT  0.930 3.760 3.140 4.000 ;
        RECT  0.930 3.760 1.170 4.610 ;
        RECT  3.690 1.610 4.260 1.850 ;
        RECT  4.020 1.610 4.260 3.380 ;
        RECT  3.690 3.140 4.260 3.380 ;
        RECT  4.980 1.620 6.100 1.860 ;
        RECT  5.860 2.170 6.310 2.570 ;
        RECT  5.860 1.620 6.100 3.720 ;
        RECT  4.980 3.480 6.100 3.720 ;
        RECT  6.340 1.610 6.880 1.930 ;
        RECT  6.640 1.610 6.880 2.840 ;
        RECT  6.670 2.600 6.910 3.720 ;
        RECT  6.340 3.480 6.910 3.720 ;
        RECT  3.030 1.130 7.360 1.370 ;
        RECT  7.120 1.130 7.360 2.340 ;
        RECT  7.230 2.100 7.470 3.450 ;
        RECT  3.030 1.130 3.270 3.460 ;
        RECT  8.530 1.770 8.920 2.090 ;
        RECT  8.530 1.770 8.770 3.450 ;
        RECT  8.530 3.130 9.060 3.450 ;
        RECT  7.780 1.770 8.230 2.090 ;
        RECT  7.990 1.770 8.230 3.930 ;
        RECT  10.580 2.520 10.820 3.930 ;
        RECT  7.990 3.690 10.820 3.930 ;
        RECT  10.100 1.850 11.300 2.090 ;
        RECT  9.010 2.380 10.340 2.620 ;
        RECT  11.060 1.850 11.300 3.370 ;
        RECT  11.060 3.130 11.860 3.370 ;
        RECT  10.100 1.850 10.340 3.450 ;
        RECT  12.210 1.850 13.260 2.090 ;
        RECT  13.020 1.850 13.260 4.160 ;
        RECT  4.500 2.520 4.740 4.200 ;
        RECT  11.210 3.920 13.890 4.160 ;
        RECT  4.500 3.960 6.580 4.200 ;
        RECT  11.210 3.920 11.450 4.410 ;
        RECT  6.340 4.170 11.450 4.410 ;
        RECT  13.650 3.920 13.890 4.570 ;
        RECT  11.540 1.370 13.740 1.610 ;
        RECT  13.500 1.540 14.510 1.780 ;
        RECT  14.270 1.540 14.510 2.250 ;
        RECT  14.270 2.010 15.120 2.250 ;
        RECT  11.540 1.370 11.780 2.890 ;
        RECT  11.540 2.650 12.520 2.890 ;
        RECT  12.280 2.650 12.520 3.450 ;
        RECT  14.750 1.480 15.600 1.720 ;
        RECT  15.360 2.010 16.080 2.250 ;
        RECT  15.050 2.610 15.600 2.850 ;
        RECT  15.360 1.480 15.600 2.850 ;
        RECT  13.500 2.850 15.290 3.090 ;
        RECT  15.050 2.610 15.290 4.220 ;
    END
END deprq1

MACRO depfq4
    CLASS CORE ;
    FOREIGN depfq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 2.580 6.100 3.020 ;
        RECT  5.660 2.100 6.030 3.020 ;
        RECT  5.630 2.100 6.030 2.500 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.385  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.740 3.020 ;
        RECT  2.300 1.950 2.660 3.020 ;
        RECT  2.250 1.950 2.660 2.350 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.990 0.880 2.390 ;
        RECT  0.120 1.990 0.500 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.960  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.540 2.580 18.920 3.020 ;
        RECT  16.470 3.620 18.900 3.860 ;
        RECT  18.600 1.510 18.900 3.860 ;
        RECT  18.570 1.190 18.810 1.750 ;
        RECT  17.000 1.510 18.900 1.750 ;
        END
    END Q
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.796  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.410 3.920 13.990 4.160 ;
        RECT  13.750 2.590 13.990 4.160 ;
        RECT  13.320 2.590 13.990 3.130 ;
        RECT  11.710 4.380 13.650 4.620 ;
        RECT  13.410 3.920 13.650 4.620 ;
        RECT  11.710 3.840 11.950 4.620 ;
        RECT  10.850 3.840 11.950 4.080 ;
        RECT  10.850 3.260 11.090 4.080 ;
        RECT  9.920 3.260 11.090 3.500 ;
        RECT  9.920 2.600 10.160 3.500 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 19.040 5.600 ;
        RECT  18.330 4.540 18.730 5.600 ;
        RECT  17.030 4.540 17.430 5.600 ;
        RECT  15.730 3.530 16.130 5.600 ;
        RECT  13.890 4.400 14.290 5.600 ;
        RECT  10.960 4.320 11.360 5.600 ;
        RECT  9.420 4.320 9.820 5.600 ;
        RECT  5.930 4.710 6.330 5.600 ;
        RECT  4.620 4.710 5.020 5.600 ;
        RECT  1.990 4.380 2.390 5.600 ;
        RECT  0.720 4.100 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 19.040 0.740 ;
        RECT  17.750 0.000 18.150 1.270 ;
        RECT  16.100 0.000 16.500 0.890 ;
        RECT  14.330 0.000 14.730 0.890 ;
        RECT  10.260 0.000 10.500 1.280 ;
        RECT  5.950 0.000 6.350 0.890 ;
        RECT  4.860 0.000 5.260 0.890 ;
        RECT  2.020 0.000 2.420 0.890 ;
        RECT  0.730 0.000 1.150 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.510 1.360 1.750 ;
        RECT  1.120 1.510 1.360 2.510 ;
        RECT  1.290 2.270 1.530 3.170 ;
        RECT  0.910 2.930 1.530 3.170 ;
        RECT  0.910 2.930 1.150 3.560 ;
        RECT  0.150 3.320 1.150 3.560 ;
        RECT  2.870 1.360 3.140 1.760 ;
        RECT  2.900 1.360 3.140 2.090 ;
        RECT  3.140 1.850 3.380 3.660 ;
        RECT  2.730 3.420 3.380 3.660 ;
        RECT  1.600 1.460 1.840 2.030 ;
        RECT  1.460 3.530 2.010 3.770 ;
        RECT  1.770 1.790 2.010 4.140 ;
        RECT  3.620 2.440 3.860 4.140 ;
        RECT  1.770 3.900 3.860 4.140 ;
        RECT  4.110 1.610 4.670 1.850 ;
        RECT  4.110 1.610 4.350 3.920 ;
        RECT  5.560 1.610 6.580 1.850 ;
        RECT  6.270 1.610 6.580 2.400 ;
        RECT  6.340 2.520 6.740 2.920 ;
        RECT  5.680 3.260 6.580 3.500 ;
        RECT  6.340 1.610 6.580 3.500 ;
        RECT  5.300 3.400 6.100 3.640 ;
        RECT  7.000 1.520 7.240 2.170 ;
        RECT  7.100 1.930 7.340 3.400 ;
        RECT  6.820 3.160 7.340 3.400 ;
        RECT  6.820 3.160 7.060 4.140 ;
        RECT  6.610 3.740 7.060 4.140 ;
        RECT  6.580 0.980 7.940 1.220 ;
        RECT  3.610 1.130 6.810 1.370 ;
        RECT  3.610 1.130 3.850 1.730 ;
        RECT  7.700 0.980 7.940 2.050 ;
        RECT  4.910 1.130 5.150 3.160 ;
        RECT  7.630 1.810 7.870 3.970 ;
        RECT  7.310 3.730 7.870 3.970 ;
        RECT  4.820 2.920 5.060 4.470 ;
        RECT  4.140 4.230 5.060 4.470 ;
        RECT  3.290 4.380 4.380 4.620 ;
        RECT  9.000 1.460 9.540 1.860 ;
        RECT  9.000 1.460 9.240 2.150 ;
        RECT  8.730 1.910 9.240 2.150 ;
        RECT  8.730 1.910 8.970 4.280 ;
        RECT  8.360 0.980 10.020 1.220 ;
        RECT  9.780 0.980 10.020 1.760 ;
        RECT  8.360 0.980 8.760 1.670 ;
        RECT  9.780 1.520 11.140 1.760 ;
        RECT  10.900 1.520 11.140 2.540 ;
        RECT  10.900 2.300 11.560 2.540 ;
        RECT  8.180 1.350 8.420 3.110 ;
        RECT  8.130 2.870 8.370 3.510 ;
        RECT  11.420 1.560 12.040 1.800 ;
        RECT  9.480 2.120 10.640 2.360 ;
        RECT  9.440 2.300 9.720 2.460 ;
        RECT  9.220 2.390 9.680 2.630 ;
        RECT  10.400 2.120 10.640 3.020 ;
        RECT  11.800 1.560 12.040 3.020 ;
        RECT  10.400 2.780 12.040 3.020 ;
        RECT  11.660 2.780 11.900 3.600 ;
        RECT  9.220 2.390 9.460 3.980 ;
        RECT  9.220 3.740 10.590 3.980 ;
        RECT  12.780 1.560 13.500 1.800 ;
        RECT  13.340 1.610 14.470 1.850 ;
        RECT  14.230 1.670 15.260 1.910 ;
        RECT  12.780 2.100 13.590 2.340 ;
        RECT  12.780 1.560 13.020 3.630 ;
        RECT  12.780 3.390 13.510 3.630 ;
        RECT  14.230 1.610 14.470 4.020 ;
        RECT  14.230 3.780 14.850 4.020 ;
        RECT  12.280 0.980 14.090 1.220 ;
        RECT  13.850 1.130 15.420 1.370 ;
        RECT  15.020 1.030 15.420 1.430 ;
        RECT  12.280 0.980 12.520 3.550 ;
        RECT  12.240 3.310 12.480 4.140 ;
        RECT  12.240 3.900 12.790 4.140 ;
        RECT  15.660 1.630 16.740 1.870 ;
        RECT  16.500 2.300 18.200 2.700 ;
        RECT  14.750 2.780 14.990 3.330 ;
        RECT  15.290 3.040 16.740 3.280 ;
        RECT  16.500 1.630 16.740 3.280 ;
        RECT  14.750 3.090 15.480 3.330 ;
        RECT  15.240 3.090 15.480 4.620 ;
    END
END depfq4

MACRO depfq2
    CLASS CORE ;
    FOREIGN depfq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.176  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.230 2.020 4.830 2.540 ;
        RECT  3.980 2.020 4.830 2.480 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.550 1.140 3.020 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.530 0.460 3.180 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.986  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.680 2.580 16.180 3.020 ;
        RECT  15.680 2.580 16.000 3.450 ;
        RECT  15.680 1.930 15.920 3.450 ;
        RECT  15.590 1.550 15.830 2.130 ;
        END
    END Q
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.940 2.300 13.610 2.700 ;
        RECT  12.940 2.300 13.380 3.020 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  16.330 3.760 16.570 5.600 ;
        RECT  15.070 4.710 15.470 5.600 ;
        RECT  13.110 4.710 13.510 5.600 ;
        RECT  9.650 4.710 10.050 5.600 ;
        RECT  8.540 4.710 8.940 5.600 ;
        RECT  5.780 4.320 6.020 5.600 ;
        RECT  4.230 4.320 4.490 5.600 ;
        RECT  3.220 4.710 3.620 5.600 ;
        RECT  0.230 3.420 1.060 3.660 ;
        RECT  0.740 3.260 1.060 3.660 ;
        RECT  0.230 3.420 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  16.330 0.000 16.570 1.550 ;
        RECT  14.850 0.000 15.090 1.620 ;
        RECT  13.520 0.000 13.920 0.890 ;
        RECT  9.800 0.000 10.200 1.040 ;
        RECT  8.180 0.000 8.580 0.890 ;
        RECT  4.330 0.000 4.730 0.890 ;
        RECT  1.830 0.000 2.230 0.900 ;
        RECT  0.230 1.780 0.820 2.020 ;
        RECT  0.230 0.000 0.470 2.020 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.860 1.700 2.100 3.600 ;
        RECT  0.930 0.980 1.600 1.220 ;
        RECT  1.310 1.210 2.510 1.450 ;
        RECT  1.310 0.980 1.550 2.380 ;
        RECT  1.380 2.210 1.620 4.610 ;
        RECT  0.890 4.370 2.100 4.610 ;
        RECT  2.340 2.670 2.580 4.400 ;
        RECT  2.750 0.980 3.680 1.220 ;
        RECT  3.340 1.720 3.580 2.910 ;
        RECT  3.560 2.670 3.800 3.600 ;
        RECT  5.220 1.610 5.460 3.520 ;
        RECT  4.840 3.270 5.460 3.520 ;
        RECT  2.520 1.720 3.060 2.040 ;
        RECT  5.720 1.770 6.360 2.090 ;
        RECT  2.820 1.720 3.060 4.080 ;
        RECT  5.720 1.770 5.960 4.080 ;
        RECT  2.820 3.840 5.960 4.080 ;
        RECT  7.330 1.760 7.850 2.050 ;
        RECT  7.330 1.760 7.570 2.540 ;
        RECT  7.220 2.300 7.460 3.550 ;
        RECT  6.670 1.770 7.090 2.090 ;
        RECT  6.670 1.770 6.910 3.070 ;
        RECT  7.700 2.890 9.540 3.130 ;
        RECT  6.480 2.820 6.720 4.030 ;
        RECT  7.700 2.890 7.940 3.990 ;
        RECT  6.480 3.790 7.910 4.030 ;
        RECT  9.490 1.760 9.730 2.630 ;
        RECT  7.810 2.390 10.020 2.630 ;
        RECT  9.780 2.390 10.020 3.730 ;
        RECT  9.670 3.340 10.060 3.730 ;
        RECT  9.780 3.260 10.060 3.730 ;
        RECT  8.700 3.490 10.060 3.730 ;
        RECT  10.570 0.980 11.640 1.220 ;
        RECT  8.080 4.230 11.510 4.470 ;
        RECT  6.520 4.380 8.310 4.620 ;
        RECT  11.240 4.380 12.150 4.620 ;
        RECT  3.970 1.130 9.220 1.370 ;
        RECT  8.990 1.280 10.210 1.520 ;
        RECT  9.970 1.280 10.210 2.040 ;
        RECT  9.970 1.800 10.540 2.040 ;
        RECT  12.350 1.770 12.590 2.850 ;
        RECT  11.600 2.610 12.590 2.850 ;
        RECT  10.300 1.800 10.540 3.930 ;
        RECT  11.600 2.610 11.840 3.930 ;
        RECT  10.300 3.690 12.370 3.930 ;
        RECT  12.120 3.890 14.080 4.130 ;
        RECT  11.870 1.290 13.260 1.530 ;
        RECT  13.020 1.290 13.260 2.060 ;
        RECT  10.860 1.770 11.410 2.090 ;
        RECT  13.020 1.820 14.100 2.060 ;
        RECT  11.870 1.290 12.110 2.090 ;
        RECT  10.860 1.850 12.110 2.090 ;
        RECT  13.860 1.820 14.100 2.840 ;
        RECT  13.860 2.600 14.680 2.840 ;
        RECT  10.860 1.770 11.100 3.450 ;
        RECT  14.030 1.300 14.600 1.540 ;
        RECT  14.360 1.300 14.600 2.160 ;
        RECT  14.360 1.920 15.330 2.160 ;
        RECT  14.380 3.110 15.330 3.360 ;
        RECT  15.090 1.920 15.330 3.360 ;
        RECT  12.750 3.300 14.780 3.540 ;
    END
END depfq2

MACRO depfq1
    CLASS CORE ;
    FOREIGN depfq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.176  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.230 2.020 4.830 2.540 ;
        RECT  3.980 2.020 4.830 2.480 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.550 1.140 3.020 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.530 0.460 3.180 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.011  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 3.700 16.210 4.140 ;
        RECT  15.970 0.980 16.210 4.140 ;
        END
    END Q
    PIN SDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.940 2.020 13.620 2.700 ;
        END
    END SDN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  15.070 4.710 15.470 5.600 ;
        RECT  13.300 4.710 13.700 5.600 ;
        RECT  9.840 4.710 10.240 5.600 ;
        RECT  8.730 4.710 9.130 5.600 ;
        RECT  5.780 4.320 6.020 5.600 ;
        RECT  4.230 4.320 4.490 5.600 ;
        RECT  3.220 4.710 3.620 5.600 ;
        RECT  0.230 3.420 1.060 3.660 ;
        RECT  0.740 3.260 1.060 3.660 ;
        RECT  0.230 3.420 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  15.000 0.000 15.400 1.050 ;
        RECT  13.520 0.000 13.920 1.050 ;
        RECT  9.800 0.000 10.200 1.040 ;
        RECT  8.180 0.000 8.580 0.890 ;
        RECT  4.330 0.000 4.730 0.890 ;
        RECT  1.830 0.000 2.230 0.900 ;
        RECT  0.230 1.780 0.820 2.020 ;
        RECT  0.230 0.000 0.470 2.020 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.860 1.700 2.100 3.600 ;
        RECT  0.930 0.980 1.600 1.220 ;
        RECT  1.310 1.210 2.510 1.450 ;
        RECT  1.310 0.980 1.550 2.380 ;
        RECT  1.380 2.210 1.620 4.610 ;
        RECT  0.890 4.370 2.100 4.610 ;
        RECT  2.340 2.670 2.580 4.400 ;
        RECT  2.750 0.980 3.680 1.220 ;
        RECT  3.340 1.720 3.580 2.910 ;
        RECT  3.560 2.670 3.800 3.600 ;
        RECT  5.220 2.670 5.670 3.070 ;
        RECT  5.220 1.610 5.460 3.520 ;
        RECT  4.840 3.270 5.460 3.520 ;
        RECT  2.520 1.720 3.060 2.040 ;
        RECT  5.940 1.770 6.430 2.090 ;
        RECT  2.820 1.720 3.060 4.080 ;
        RECT  5.940 1.770 6.180 4.080 ;
        RECT  2.820 3.840 6.180 4.080 ;
        RECT  7.520 1.760 7.920 2.050 ;
        RECT  7.520 1.760 7.760 3.550 ;
        RECT  6.700 1.770 7.160 2.090 ;
        RECT  8.560 2.890 9.720 3.130 ;
        RECT  8.560 2.890 8.800 3.600 ;
        RECT  8.080 3.360 8.800 3.600 ;
        RECT  6.700 1.770 6.940 4.030 ;
        RECT  7.930 3.750 8.320 3.990 ;
        RECT  8.080 3.360 8.320 3.990 ;
        RECT  6.700 3.790 8.130 4.030 ;
        RECT  9.490 1.760 9.730 2.520 ;
        RECT  8.000 2.280 10.200 2.520 ;
        RECT  8.000 2.280 8.400 2.710 ;
        RECT  9.960 2.280 10.200 3.730 ;
        RECT  9.960 3.270 10.270 3.730 ;
        RECT  9.040 3.370 10.270 3.730 ;
        RECT  10.570 0.980 11.640 1.220 ;
        RECT  8.270 4.230 12.340 4.470 ;
        RECT  6.520 4.380 8.500 4.620 ;
        RECT  3.970 1.130 9.220 1.370 ;
        RECT  8.990 1.280 10.210 1.520 ;
        RECT  9.970 1.280 10.210 2.040 ;
        RECT  9.970 1.800 10.750 2.040 ;
        RECT  12.350 1.770 12.590 2.850 ;
        RECT  11.810 2.610 12.590 2.850 ;
        RECT  10.510 1.800 10.750 3.930 ;
        RECT  11.810 2.610 12.050 3.930 ;
        RECT  10.510 3.690 14.290 3.930 ;
        RECT  11.870 1.290 14.100 1.530 ;
        RECT  10.990 1.770 11.410 2.090 ;
        RECT  11.870 1.290 12.110 2.090 ;
        RECT  10.990 1.850 12.110 2.090 ;
        RECT  10.990 1.770 11.310 2.170 ;
        RECT  13.860 1.290 14.100 2.840 ;
        RECT  13.860 2.600 15.150 2.840 ;
        RECT  11.070 1.770 11.310 3.450 ;
        RECT  14.340 0.980 14.580 1.530 ;
        RECT  14.340 1.290 15.630 1.530 ;
        RECT  15.390 1.290 15.630 3.340 ;
        RECT  12.760 3.100 15.630 3.340 ;
        RECT  14.590 3.100 14.990 3.450 ;
    END
END depfq1

MACRO denrq4
    CLASS CORE ;
    FOREIGN denrq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.560 2.460 6.960 2.860 ;
        RECT  6.220 2.580 6.660 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.290 2.580 2.740 3.020 ;
        RECT  2.290 2.330 2.710 3.020 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.320 0.780 2.720 ;
        RECT  0.120 2.320 0.500 3.020 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.893  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.420 2.440 17.800 3.020 ;
        RECT  17.200 1.250 17.440 2.680 ;
        RECT  15.220 2.440 17.800 2.680 ;
        RECT  17.030 1.250 17.440 1.650 ;
        RECT  15.660 1.350 17.440 1.590 ;
        RECT  16.420 2.440 16.660 4.320 ;
        RECT  15.220 2.440 15.620 2.950 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 17.920 5.600 ;
        RECT  17.050 4.120 17.450 5.600 ;
        RECT  15.780 3.230 16.180 5.600 ;
        RECT  14.440 4.470 14.840 5.600 ;
        RECT  10.890 4.710 11.290 5.600 ;
        RECT  7.490 4.690 7.890 5.600 ;
        RECT  6.310 4.690 6.710 5.600 ;
        RECT  4.850 4.690 5.250 5.600 ;
        RECT  2.160 4.110 2.560 5.600 ;
        RECT  0.800 4.160 1.200 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 17.920 0.740 ;
        RECT  16.240 0.000 16.640 0.980 ;
        RECT  14.870 0.000 15.270 0.890 ;
        RECT  14.130 0.000 14.530 0.890 ;
        RECT  10.590 0.000 10.990 0.890 ;
        RECT  6.970 0.000 7.370 1.090 ;
        RECT  4.910 0.000 5.310 1.160 ;
        RECT  2.210 0.000 2.610 0.980 ;
        RECT  0.740 0.000 1.140 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.780 1.260 2.020 ;
        RECT  1.020 2.270 1.540 2.670 ;
        RECT  1.020 1.780 1.260 3.550 ;
        RECT  0.150 3.310 1.260 3.550 ;
        RECT  2.800 1.780 3.420 2.020 ;
        RECT  3.180 1.780 3.420 3.010 ;
        RECT  2.980 2.770 3.220 3.830 ;
        RECT  2.730 3.430 3.220 3.830 ;
        RECT  3.730 1.040 4.470 1.280 ;
        RECT  1.510 1.220 3.970 1.460 ;
        RECT  1.510 1.220 2.020 1.900 ;
        RECT  1.780 1.220 2.020 3.150 ;
        RECT  1.540 2.910 1.780 3.500 ;
        RECT  4.140 1.780 4.720 2.020 ;
        RECT  4.140 1.780 4.380 3.490 ;
        RECT  4.150 3.220 4.650 3.620 ;
        RECT  5.630 1.690 6.080 2.090 ;
        RECT  4.620 2.500 5.870 2.740 ;
        RECT  5.630 1.690 5.870 3.620 ;
        RECT  6.380 1.510 7.440 1.750 ;
        RECT  7.200 2.230 7.880 2.470 ;
        RECT  7.200 1.510 7.440 3.610 ;
        RECT  6.900 3.210 7.440 3.610 ;
        RECT  8.600 1.610 8.840 2.400 ;
        RECT  8.600 2.160 9.360 2.400 ;
        RECT  3.660 1.700 3.900 4.100 ;
        RECT  3.510 3.590 3.910 4.100 ;
        RECT  3.510 3.860 9.360 4.100 ;
        RECT  9.120 2.160 9.360 4.130 ;
        RECT  8.900 3.730 9.360 4.130 ;
        RECT  10.080 1.610 10.320 3.380 ;
        RECT  10.080 3.140 10.660 3.380 ;
        RECT  9.260 1.580 9.840 1.820 ;
        RECT  11.080 2.610 11.700 2.850 ;
        RECT  9.600 1.580 9.840 3.860 ;
        RECT  11.080 2.610 11.320 3.860 ;
        RECT  9.600 3.620 11.320 3.860 ;
        RECT  7.740 0.980 10.280 1.220 ;
        RECT  11.430 1.020 12.210 1.260 ;
        RECT  10.030 1.130 11.670 1.370 ;
        RECT  7.740 0.980 8.360 1.800 ;
        RECT  8.120 0.980 8.360 3.580 ;
        RECT  8.120 2.640 8.790 3.040 ;
        RECT  8.120 2.640 8.600 3.580 ;
        RECT  11.190 1.620 11.850 1.860 ;
        RECT  11.190 1.620 11.430 2.370 ;
        RECT  10.580 2.130 12.260 2.370 ;
        RECT  10.580 2.130 10.820 2.740 ;
        RECT  12.020 2.130 12.260 3.380 ;
        RECT  11.660 3.140 12.260 3.380 ;
        RECT  10.170 4.230 11.930 4.470 ;
        RECT  11.690 4.290 12.420 4.530 ;
        RECT  8.730 4.380 10.410 4.620 ;
        RECT  13.010 1.580 13.250 3.460 ;
        RECT  13.010 3.060 13.570 3.460 ;
        RECT  13.270 3.060 13.510 4.610 ;
        RECT  12.510 1.000 13.860 1.240 ;
        RECT  12.190 1.630 12.750 1.870 ;
        RECT  13.620 1.000 13.860 2.140 ;
        RECT  13.620 1.900 14.400 2.140 ;
        RECT  12.510 1.000 12.750 3.460 ;
        RECT  14.320 1.350 14.880 1.590 ;
        RECT  14.640 1.940 16.960 2.180 ;
        RECT  14.640 1.350 14.880 3.860 ;
        RECT  13.870 3.620 14.880 3.860 ;
    END
END denrq4

MACRO denrq2
    CLASS CORE ;
    FOREIGN denrq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.178  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.580 5.990 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.086  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.700 2.740 4.590 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.580 2.700 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.050 2.580 15.620 3.020 ;
        RECT  15.050 1.690 15.290 3.460 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  15.700 4.080 15.940 5.600 ;
        RECT  14.390 4.080 14.630 5.600 ;
        RECT  12.700 4.710 13.100 5.600 ;
        RECT  9.810 4.710 10.210 5.600 ;
        RECT  5.930 4.710 6.330 5.600 ;
        RECT  4.640 4.710 5.040 5.600 ;
        RECT  1.690 4.710 2.090 5.600 ;
        RECT  0.970 4.430 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  15.740 0.000 15.980 1.400 ;
        RECT  14.190 0.000 14.430 1.460 ;
        RECT  12.650 0.000 13.050 0.890 ;
        RECT  9.860 0.000 10.100 1.930 ;
        RECT  5.930 0.000 6.330 0.890 ;
        RECT  4.640 0.000 5.040 0.890 ;
        RECT  1.620 0.000 2.020 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 2.460 1.570 2.700 ;
        RECT  0.820 1.770 1.060 3.180 ;
        RECT  0.230 2.940 1.060 3.180 ;
        RECT  0.230 2.940 0.470 4.600 ;
        RECT  2.410 1.610 2.650 3.460 ;
        RECT  0.850 1.040 1.250 1.370 ;
        RECT  0.850 1.130 3.150 1.370 ;
        RECT  2.910 1.130 3.150 2.910 ;
        RECT  1.820 1.130 2.060 3.660 ;
        RECT  0.920 3.420 2.060 3.660 ;
        RECT  4.130 1.610 4.370 3.720 ;
        RECT  5.340 1.690 6.470 1.930 ;
        RECT  6.230 2.170 6.670 2.570 ;
        RECT  6.230 1.690 6.470 3.910 ;
        RECT  5.340 3.670 6.470 3.910 ;
        RECT  6.710 1.610 7.210 1.930 ;
        RECT  6.970 1.610 7.210 3.990 ;
        RECT  6.710 3.670 7.210 3.990 ;
        RECT  3.390 1.130 7.740 1.370 ;
        RECT  7.500 1.130 7.740 3.510 ;
        RECT  3.390 1.130 3.630 3.720 ;
        RECT  9.120 1.770 9.360 3.510 ;
        RECT  9.600 2.900 10.680 3.140 ;
        RECT  8.240 1.770 8.480 3.990 ;
        RECT  9.600 2.900 9.840 3.990 ;
        RECT  8.240 3.750 9.840 3.990 ;
        RECT  10.610 1.770 10.850 2.620 ;
        RECT  9.600 2.380 11.160 2.620 ;
        RECT  10.920 2.380 11.160 3.670 ;
        RECT  10.560 3.430 11.160 3.670 ;
        RECT  4.290 3.960 4.700 4.470 ;
        RECT  12.140 1.710 12.380 4.470 ;
        RECT  4.290 4.230 12.380 4.470 ;
        RECT  11.400 1.230 13.310 1.470 ;
        RECT  13.070 1.230 13.310 2.700 ;
        RECT  11.400 1.230 11.640 3.750 ;
        RECT  13.550 1.690 13.790 3.460 ;
        RECT  13.550 2.390 14.810 2.630 ;
        RECT  12.670 3.060 13.820 3.300 ;
        RECT  13.550 2.390 13.820 3.460 ;
        RECT  13.420 3.060 13.820 3.460 ;
    END
END denrq2

MACRO denrq1
    CLASS CORE ;
    FOREIGN denrq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.178  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.580 5.990 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.086  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.700 2.740 4.590 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.580 2.700 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.620 3.060 15.370 3.580 ;
        RECT  15.050 1.690 15.370 3.580 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.680 5.600 ;
        RECT  14.390 4.080 14.630 5.600 ;
        RECT  12.700 4.710 13.100 5.600 ;
        RECT  9.810 4.710 10.210 5.600 ;
        RECT  5.930 4.710 6.330 5.600 ;
        RECT  4.640 4.710 5.040 5.600 ;
        RECT  1.690 4.710 2.090 5.600 ;
        RECT  0.970 4.430 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.680 0.740 ;
        RECT  14.190 0.000 14.430 1.460 ;
        RECT  12.650 0.000 13.050 0.890 ;
        RECT  9.860 0.000 10.100 1.930 ;
        RECT  5.930 0.000 6.330 0.890 ;
        RECT  4.640 0.000 5.040 0.890 ;
        RECT  1.620 0.000 2.020 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 2.460 1.570 2.700 ;
        RECT  0.820 1.770 1.060 3.180 ;
        RECT  0.230 2.940 1.060 3.180 ;
        RECT  0.230 2.940 0.470 4.600 ;
        RECT  2.410 1.610 2.650 3.460 ;
        RECT  0.850 1.040 1.250 1.370 ;
        RECT  0.850 1.130 3.150 1.370 ;
        RECT  2.910 1.130 3.150 2.910 ;
        RECT  1.820 1.130 2.060 3.660 ;
        RECT  0.920 3.420 2.060 3.660 ;
        RECT  4.130 1.610 4.370 3.720 ;
        RECT  5.340 1.690 6.470 1.930 ;
        RECT  6.230 2.170 6.670 2.570 ;
        RECT  6.230 1.690 6.470 3.910 ;
        RECT  5.340 3.670 6.470 3.910 ;
        RECT  6.710 1.610 7.210 1.930 ;
        RECT  6.970 1.610 7.210 3.990 ;
        RECT  6.710 3.670 7.210 3.990 ;
        RECT  3.390 1.130 7.740 1.370 ;
        RECT  7.500 1.130 7.740 3.510 ;
        RECT  3.390 1.130 3.630 3.720 ;
        RECT  9.120 1.770 9.360 3.510 ;
        RECT  9.600 2.900 10.680 3.140 ;
        RECT  8.240 1.770 8.480 3.990 ;
        RECT  9.600 2.900 9.840 3.990 ;
        RECT  8.240 3.750 9.840 3.990 ;
        RECT  10.610 1.770 10.850 2.620 ;
        RECT  9.600 2.380 11.160 2.620 ;
        RECT  10.920 2.380 11.160 3.670 ;
        RECT  10.560 3.430 11.160 3.670 ;
        RECT  4.290 3.960 4.700 4.470 ;
        RECT  12.140 1.710 12.380 4.470 ;
        RECT  4.290 4.230 12.380 4.470 ;
        RECT  11.400 1.230 13.310 1.470 ;
        RECT  13.070 1.230 13.310 2.700 ;
        RECT  11.400 1.230 11.640 3.750 ;
        RECT  13.550 1.690 13.790 3.460 ;
        RECT  13.550 2.300 14.810 2.540 ;
        RECT  12.670 3.060 13.820 3.300 ;
        RECT  13.550 2.300 13.820 3.460 ;
        RECT  13.420 3.060 13.820 3.460 ;
    END
END denrq1

MACRO decrq4
    CLASS CORE ;
    FOREIGN decrq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.875  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.020 4.070 16.530 4.310 ;
        RECT  16.290 2.430 16.530 4.310 ;
        RECT  13.790 3.860 15.260 4.100 ;
        RECT  12.190 4.380 14.030 4.620 ;
        RECT  13.790 3.860 14.030 4.620 ;
        RECT  12.190 3.690 12.430 4.620 ;
        RECT  11.440 3.690 12.430 3.930 ;
        RECT  11.440 2.580 11.700 3.930 ;
        RECT  11.220 2.110 11.460 3.160 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.800 2.780 6.660 3.020 ;
        RECT  6.160 2.580 6.660 3.020 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 1.910 2.780 2.460 ;
        RECT  2.350 1.910 2.590 2.880 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.380 0.980 2.620 ;
        RECT  0.120 2.380 0.500 3.030 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.497  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.840 3.520 20.600 3.920 ;
        RECT  20.150 1.370 20.600 3.920 ;
        RECT  18.190 1.370 20.600 1.770 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.720 5.600 ;
        RECT  19.900 4.320 20.300 5.600 ;
        RECT  18.600 4.320 19.000 5.600 ;
        RECT  17.230 4.180 17.630 5.600 ;
        RECT  16.430 4.650 16.830 5.600 ;
        RECT  15.030 4.690 15.430 5.600 ;
        RECT  14.310 4.340 14.550 5.600 ;
        RECT  11.430 4.710 11.830 5.600 ;
        RECT  9.950 4.710 10.350 5.600 ;
        RECT  5.700 4.710 6.100 5.600 ;
        RECT  5.000 4.710 5.400 5.600 ;
        RECT  2.210 4.570 2.610 5.600 ;
        RECT  0.760 4.330 1.160 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.720 0.740 ;
        RECT  18.980 0.000 19.380 1.100 ;
        RECT  17.450 0.000 17.850 1.210 ;
        RECT  16.480 0.000 16.720 1.160 ;
        RECT  14.350 0.000 14.750 0.890 ;
        RECT  11.310 0.000 11.710 0.890 ;
        RECT  7.160 0.000 7.560 0.890 ;
        RECT  5.690 0.000 5.930 1.660 ;
        RECT  1.970 0.000 2.370 0.890 ;
        RECT  1.020 0.000 1.420 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 0.980 0.460 2.090 ;
        RECT  0.180 1.480 0.590 2.090 ;
        RECT  0.180 1.850 1.460 2.090 ;
        RECT  1.220 1.850 1.460 3.510 ;
        RECT  0.260 3.270 1.460 3.510 ;
        RECT  0.260 3.270 0.500 3.900 ;
        RECT  3.040 1.560 3.280 2.360 ;
        RECT  3.020 2.120 3.260 3.490 ;
        RECT  2.780 3.090 3.260 3.490 ;
        RECT  2.620 0.980 4.570 1.220 ;
        RECT  1.770 1.160 2.860 1.400 ;
        RECT  4.330 0.980 4.570 1.830 ;
        RECT  4.460 1.600 4.700 2.250 ;
        RECT  4.460 1.840 4.940 2.250 ;
        RECT  1.770 1.160 2.010 3.520 ;
        RECT  1.820 3.280 2.060 4.030 ;
        RECT  1.820 3.740 3.740 3.980 ;
        RECT  3.500 2.520 3.740 3.980 ;
        RECT  1.510 3.790 2.630 4.030 ;
        RECT  4.870 1.190 5.440 1.430 ;
        RECT  5.200 1.190 5.440 2.740 ;
        RECT  4.460 2.500 5.440 2.740 ;
        RECT  4.460 2.500 4.700 3.550 ;
        RECT  6.190 0.980 6.920 1.220 ;
        RECT  6.680 0.980 6.920 1.870 ;
        RECT  6.360 1.630 7.140 1.870 ;
        RECT  6.410 3.260 7.140 3.500 ;
        RECT  6.900 1.630 7.140 3.500 ;
        RECT  5.730 3.470 6.650 3.710 ;
        RECT  8.630 1.460 8.870 2.190 ;
        RECT  7.960 1.950 8.870 2.190 ;
        RECT  3.850 1.540 4.090 2.300 ;
        RECT  3.980 2.060 4.220 4.460 ;
        RECT  3.590 4.220 6.640 4.460 ;
        RECT  7.960 1.950 8.200 4.620 ;
        RECT  6.400 4.380 8.200 4.620 ;
        RECT  10.160 1.460 10.400 2.250 ;
        RECT  9.590 2.010 10.400 2.250 ;
        RECT  9.590 2.010 9.830 3.150 ;
        RECT  9.310 2.910 9.830 3.150 ;
        RECT  9.310 2.910 9.550 3.990 ;
        RECT  9.310 3.750 10.970 3.990 ;
        RECT  9.110 1.530 9.690 1.770 ;
        RECT  9.110 1.530 9.350 2.670 ;
        RECT  8.710 2.430 9.350 2.670 ;
        RECT  8.710 2.430 8.950 4.470 ;
        RECT  8.710 4.230 11.510 4.470 ;
        RECT  10.710 1.620 12.650 1.860 ;
        RECT  12.410 1.620 12.650 2.640 ;
        RECT  12.030 2.400 12.650 2.640 ;
        RECT  10.710 1.620 10.950 2.830 ;
        RECT  10.070 2.590 10.950 2.830 ;
        RECT  12.030 2.400 12.270 3.430 ;
        RECT  12.030 3.190 12.650 3.430 ;
        RECT  7.830 0.980 11.080 1.220 ;
        RECT  11.940 0.980 13.010 1.220 ;
        RECT  10.840 1.140 12.180 1.380 ;
        RECT  7.830 0.980 8.150 1.710 ;
        RECT  7.380 1.310 8.150 1.710 ;
        RECT  7.380 1.310 7.620 4.140 ;
        RECT  7.060 3.900 7.620 4.140 ;
        RECT  12.940 1.470 13.180 3.580 ;
        RECT  15.270 2.430 15.510 3.580 ;
        RECT  12.940 3.340 15.510 3.580 ;
        RECT  13.210 3.340 13.450 4.060 ;
        RECT  12.830 3.820 13.450 4.060 ;
        RECT  15.040 1.010 16.230 1.250 ;
        RECT  13.960 1.130 15.280 1.370 ;
        RECT  15.990 1.010 16.230 1.710 ;
        RECT  15.990 1.470 17.330 1.710 ;
        RECT  13.960 1.130 14.200 1.810 ;
        RECT  13.420 1.570 14.200 1.810 ;
        RECT  13.420 1.570 13.660 3.100 ;
        RECT  13.420 2.860 14.010 3.100 ;
        RECT  14.720 1.630 15.730 1.870 ;
        RECT  15.490 1.630 15.730 2.190 ;
        RECT  15.490 1.950 17.540 2.190 ;
        RECT  14.720 1.630 14.960 2.350 ;
        RECT  14.070 2.110 14.960 2.350 ;
        RECT  17.300 2.040 19.810 2.460 ;
        RECT  15.790 1.950 16.030 3.610 ;
    END
END decrq4

MACRO decrq2
    CLASS CORE ;
    FOREIGN decrq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.500 3.140 14.240 3.580 ;
        RECT  13.840 2.930 14.240 3.580 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.218  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 3.140 4.980 3.580 ;
        RECT  4.540 2.520 4.850 3.580 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.169  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.370 1.010 3.020 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 1.900 ;
        RECT  0.120 3.260 0.460 3.660 ;
        RECT  0.120 1.460 0.360 3.660 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.377  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.180 2.020 15.620 3.480 ;
        RECT  15.180 1.100 15.420 3.480 ;
        RECT  14.940 1.100 15.420 1.500 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  15.750 4.090 15.990 5.600 ;
        RECT  14.420 4.300 14.660 5.600 ;
        RECT  12.780 4.300 13.020 5.600 ;
        RECT  8.290 4.570 8.690 5.600 ;
        RECT  7.360 4.710 7.760 5.600 ;
        RECT  4.220 4.460 4.460 5.600 ;
        RECT  2.930 4.670 3.330 5.600 ;
        RECT  0.230 3.900 1.010 4.140 ;
        RECT  0.770 3.260 1.010 4.140 ;
        RECT  0.230 3.900 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  15.760 0.000 16.000 1.540 ;
        RECT  14.280 0.000 14.520 1.500 ;
        RECT  12.050 0.000 12.450 1.010 ;
        RECT  8.590 0.000 8.990 0.890 ;
        RECT  4.190 0.000 4.590 0.890 ;
        RECT  2.080 0.000 2.490 0.890 ;
        RECT  0.770 0.000 1.010 2.130 ;
        RECT  0.150 0.000 1.010 1.140 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.730 1.730 1.970 3.560 ;
        RECT  1.250 0.980 1.620 1.490 ;
        RECT  1.250 1.250 2.150 1.490 ;
        RECT  1.250 0.980 1.490 4.620 ;
        RECT  0.890 4.380 1.820 4.620 ;
        RECT  2.210 2.630 2.460 4.480 ;
        RECT  3.450 1.730 3.690 3.740 ;
        RECT  2.860 0.980 3.440 1.220 ;
        RECT  3.200 0.980 3.440 1.490 ;
        RECT  3.200 1.250 3.800 1.490 ;
        RECT  4.960 1.730 5.420 2.050 ;
        RECT  5.180 1.730 5.420 2.800 ;
        RECT  5.180 2.400 5.640 2.800 ;
        RECT  5.220 2.400 5.460 3.450 ;
        RECT  5.660 1.520 6.120 1.840 ;
        RECT  5.880 1.520 6.120 3.450 ;
        RECT  5.720 3.050 6.340 3.450 ;
        RECT  2.710 1.730 2.950 4.220 ;
        RECT  5.720 3.050 5.960 4.220 ;
        RECT  2.710 3.980 5.960 4.220 ;
        RECT  7.140 1.520 7.510 1.840 ;
        RECT  7.270 1.520 7.510 3.330 ;
        RECT  7.270 3.090 9.180 3.330 ;
        RECT  6.480 1.520 6.720 2.440 ;
        RECT  6.480 2.200 7.000 2.440 ;
        RECT  6.760 2.200 7.000 3.810 ;
        RECT  6.760 3.570 9.140 3.810 ;
        RECT  8.900 3.610 9.570 3.850 ;
        RECT  9.260 1.730 9.500 2.600 ;
        RECT  8.160 2.050 8.400 2.600 ;
        RECT  9.260 2.340 10.050 2.600 ;
        RECT  8.160 2.360 10.050 2.600 ;
        RECT  9.810 2.340 10.050 3.660 ;
        RECT  10.220 0.980 11.070 1.220 ;
        RECT  10.220 0.980 10.460 1.530 ;
        RECT  6.200 3.840 6.520 4.290 ;
        RECT  6.200 4.050 8.440 4.290 ;
        RECT  8.200 4.090 9.580 4.330 ;
        RECT  9.340 4.090 9.580 4.620 ;
        RECT  9.340 4.380 11.580 4.620 ;
        RECT  5.050 1.040 8.400 1.280 ;
        RECT  4.260 1.160 5.290 1.400 ;
        RECT  8.160 1.200 9.980 1.440 ;
        RECT  9.740 1.200 9.980 2.100 ;
        RECT  9.740 1.860 10.530 2.100 ;
        RECT  4.260 1.160 4.500 2.120 ;
        RECT  3.930 1.880 4.500 2.120 ;
        RECT  3.930 1.880 4.170 2.660 ;
        RECT  11.790 1.730 12.030 2.740 ;
        RECT  11.510 2.500 12.030 2.740 ;
        RECT  11.510 3.600 12.630 3.840 ;
        RECT  10.290 1.860 10.530 4.140 ;
        RECT  11.510 2.500 11.750 4.140 ;
        RECT  10.290 3.900 11.750 4.140 ;
        RECT  11.310 1.250 12.840 1.490 ;
        RECT  11.310 1.250 11.550 2.050 ;
        RECT  10.770 1.730 11.550 2.050 ;
        RECT  12.600 1.250 12.840 2.580 ;
        RECT  12.600 2.340 13.650 2.580 ;
        RECT  10.770 1.730 11.010 3.660 ;
        RECT  13.080 1.370 13.320 1.980 ;
        RECT  13.080 1.740 14.940 1.980 ;
        RECT  12.470 3.010 13.110 3.250 ;
        RECT  12.870 3.010 13.110 4.060 ;
        RECT  14.700 1.740 14.940 4.060 ;
        RECT  12.870 3.820 14.940 4.060 ;
    END
END decrq2

MACRO decrq1
    CLASS CORE ;
    FOREIGN decrq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.500 3.140 14.390 3.580 ;
        RECT  13.990 2.930 14.390 3.580 ;
        END
    END CDN
    PIN CP
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.218  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 3.140 4.980 3.580 ;
        RECT  4.540 2.520 4.850 3.580 ;
        END
    END CP
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.169  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.370 1.010 3.020 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 1.900 ;
        RECT  0.120 3.260 0.460 3.660 ;
        RECT  0.120 1.460 0.360 3.660 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.295  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.180 1.460 15.560 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.680 5.600 ;
        RECT  14.420 4.300 14.660 5.600 ;
        RECT  12.530 4.320 12.770 5.600 ;
        RECT  8.290 4.570 8.690 5.600 ;
        RECT  7.360 4.710 7.760 5.600 ;
        RECT  4.220 4.460 4.460 5.600 ;
        RECT  2.930 4.670 3.330 5.600 ;
        RECT  0.230 3.900 1.010 4.140 ;
        RECT  0.770 3.260 1.010 4.140 ;
        RECT  0.230 3.900 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.680 0.740 ;
        RECT  14.380 0.000 14.620 1.500 ;
        RECT  12.150 0.000 12.550 1.010 ;
        RECT  8.690 0.000 9.090 0.890 ;
        RECT  4.190 0.000 4.590 0.890 ;
        RECT  2.080 0.000 2.490 0.890 ;
        RECT  0.770 0.000 1.010 2.130 ;
        RECT  0.150 0.000 1.010 1.140 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.730 1.730 1.970 3.560 ;
        RECT  1.250 0.980 1.620 1.490 ;
        RECT  1.250 1.250 2.150 1.490 ;
        RECT  1.250 0.980 1.490 4.620 ;
        RECT  0.890 4.380 1.820 4.620 ;
        RECT  2.210 2.630 2.460 4.480 ;
        RECT  3.450 1.730 3.690 3.740 ;
        RECT  2.860 0.980 3.440 1.220 ;
        RECT  3.200 0.980 3.440 1.490 ;
        RECT  3.200 1.250 3.800 1.490 ;
        RECT  4.960 1.730 5.330 2.050 ;
        RECT  5.090 1.730 5.330 2.840 ;
        RECT  5.090 2.440 5.640 2.840 ;
        RECT  5.220 2.440 5.460 3.450 ;
        RECT  5.660 1.730 6.120 2.050 ;
        RECT  5.880 1.730 6.120 3.450 ;
        RECT  5.760 3.050 6.340 3.450 ;
        RECT  2.710 1.730 2.950 4.220 ;
        RECT  5.760 3.050 6.000 4.220 ;
        RECT  2.710 3.980 6.000 4.220 ;
        RECT  7.140 1.810 7.970 2.050 ;
        RECT  7.730 1.810 7.970 3.330 ;
        RECT  7.420 3.090 9.180 3.330 ;
        RECT  6.400 1.730 6.820 2.050 ;
        RECT  6.580 1.730 6.820 3.450 ;
        RECT  6.580 3.050 7.180 3.450 ;
        RECT  6.940 3.050 7.180 3.810 ;
        RECT  6.940 3.570 9.140 3.810 ;
        RECT  8.900 3.610 9.570 3.850 ;
        RECT  9.360 1.730 9.600 2.580 ;
        RECT  8.350 2.340 10.050 2.580 ;
        RECT  9.810 2.340 10.050 3.660 ;
        RECT  10.320 0.980 11.170 1.220 ;
        RECT  10.320 0.980 10.560 1.530 ;
        RECT  6.240 3.840 6.560 4.290 ;
        RECT  6.240 4.050 8.440 4.290 ;
        RECT  8.200 4.090 9.580 4.330 ;
        RECT  9.340 4.090 9.580 4.620 ;
        RECT  9.340 4.380 11.390 4.620 ;
        RECT  4.260 1.250 10.080 1.490 ;
        RECT  9.840 1.250 10.080 2.100 ;
        RECT  9.840 1.860 10.530 2.100 ;
        RECT  4.260 1.250 4.500 2.120 ;
        RECT  3.930 1.880 4.500 2.120 ;
        RECT  3.930 1.880 4.170 2.660 ;
        RECT  11.890 1.730 12.130 2.740 ;
        RECT  11.510 2.500 12.130 2.740 ;
        RECT  11.510 3.600 12.630 3.840 ;
        RECT  10.290 1.860 10.530 4.140 ;
        RECT  11.510 2.500 11.750 4.140 ;
        RECT  10.290 3.900 11.750 4.140 ;
        RECT  11.410 1.250 12.840 1.490 ;
        RECT  11.410 1.250 11.650 2.050 ;
        RECT  10.770 1.810 11.650 2.050 ;
        RECT  12.600 1.250 12.840 2.580 ;
        RECT  12.600 2.340 13.700 2.580 ;
        RECT  10.770 1.810 11.010 3.660 ;
        RECT  13.180 1.370 13.420 1.980 ;
        RECT  13.180 1.740 14.940 1.980 ;
        RECT  12.470 3.010 13.110 3.250 ;
        RECT  12.870 3.010 13.110 4.060 ;
        RECT  14.700 1.740 14.940 4.060 ;
        RECT  12.870 3.820 14.940 4.060 ;
    END
END decrq1

MACRO decfq4
    CLASS CORE ;
    FOREIGN decfq4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.872  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.020 4.070 16.530 4.310 ;
        RECT  16.290 2.430 16.530 4.310 ;
        RECT  13.790 3.860 15.260 4.100 ;
        RECT  12.190 4.380 14.030 4.620 ;
        RECT  13.790 3.860 14.030 4.620 ;
        RECT  12.190 3.690 12.430 4.620 ;
        RECT  11.440 3.690 12.430 3.930 ;
        RECT  11.440 2.580 11.700 3.930 ;
        RECT  11.220 2.120 11.460 3.160 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.493  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.800 2.780 6.660 3.020 ;
        RECT  6.160 2.580 6.660 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 2.020 2.780 2.460 ;
        RECT  2.350 2.020 2.590 2.890 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.380 0.980 2.620 ;
        RECT  0.120 2.380 0.500 3.030 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.372  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.840 3.520 20.600 3.920 ;
        RECT  20.150 1.370 20.600 3.920 ;
        RECT  18.190 1.370 20.600 1.770 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.720 5.600 ;
        RECT  19.930 4.320 20.330 5.600 ;
        RECT  18.590 4.310 18.990 5.600 ;
        RECT  17.230 4.180 17.630 5.600 ;
        RECT  16.430 4.650 16.830 5.600 ;
        RECT  15.030 4.690 15.430 5.600 ;
        RECT  14.310 4.340 14.550 5.600 ;
        RECT  11.430 4.710 11.830 5.600 ;
        RECT  9.950 4.710 10.350 5.600 ;
        RECT  5.700 4.710 6.100 5.600 ;
        RECT  5.000 4.710 5.400 5.600 ;
        RECT  2.210 4.360 2.610 5.600 ;
        RECT  0.760 4.330 1.160 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.720 0.740 ;
        RECT  18.980 0.000 19.380 1.120 ;
        RECT  17.530 0.000 17.770 1.250 ;
        RECT  16.480 0.000 16.720 1.140 ;
        RECT  14.350 0.000 14.750 0.890 ;
        RECT  11.310 0.000 11.710 0.890 ;
        RECT  7.160 0.000 7.560 0.890 ;
        RECT  5.690 0.000 5.930 1.660 ;
        RECT  1.990 0.000 2.390 0.890 ;
        RECT  1.020 0.000 1.420 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.980 0.580 2.090 ;
        RECT  0.180 1.850 1.460 2.090 ;
        RECT  1.220 1.850 1.460 3.510 ;
        RECT  0.260 3.270 1.460 3.510 ;
        RECT  0.260 3.270 0.500 3.900 ;
        RECT  3.040 1.560 3.280 2.360 ;
        RECT  3.020 2.120 3.260 3.500 ;
        RECT  2.760 3.090 3.260 3.500 ;
        RECT  2.620 0.980 4.570 1.220 ;
        RECT  1.770 1.160 2.860 1.400 ;
        RECT  4.330 0.980 4.570 1.830 ;
        RECT  4.460 1.600 4.700 2.240 ;
        RECT  4.460 1.840 4.960 2.240 ;
        RECT  1.770 1.160 2.010 4.120 ;
        RECT  3.130 3.740 3.740 3.980 ;
        RECT  3.500 2.520 3.740 3.980 ;
        RECT  1.510 3.880 3.370 4.120 ;
        RECT  1.510 3.800 1.920 4.200 ;
        RECT  4.870 1.190 5.440 1.430 ;
        RECT  5.200 1.190 5.440 2.770 ;
        RECT  4.460 2.530 5.440 2.770 ;
        RECT  4.460 2.530 4.700 3.510 ;
        RECT  6.190 0.980 6.920 1.220 ;
        RECT  6.680 0.980 6.920 1.870 ;
        RECT  6.370 1.630 7.140 1.870 ;
        RECT  6.410 3.260 7.140 3.500 ;
        RECT  6.900 1.630 7.140 3.500 ;
        RECT  5.730 3.470 6.650 3.710 ;
        RECT  8.630 1.460 8.870 2.180 ;
        RECT  8.230 1.940 8.870 2.180 ;
        RECT  3.850 1.540 4.090 2.300 ;
        RECT  8.230 1.940 8.470 3.290 ;
        RECT  7.960 3.050 8.470 3.290 ;
        RECT  3.980 2.060 4.220 4.470 ;
        RECT  3.590 4.220 4.220 4.460 ;
        RECT  3.980 4.230 6.690 4.470 ;
        RECT  7.960 3.050 8.200 4.620 ;
        RECT  6.450 4.380 8.200 4.620 ;
        RECT  10.160 1.460 10.400 2.250 ;
        RECT  9.590 2.010 10.400 2.250 ;
        RECT  9.590 2.010 9.830 3.140 ;
        RECT  9.310 2.900 9.830 3.140 ;
        RECT  9.310 2.900 9.550 3.990 ;
        RECT  9.310 3.750 10.970 3.990 ;
        RECT  9.110 1.530 9.720 1.770 ;
        RECT  9.110 1.530 9.350 2.660 ;
        RECT  8.710 2.420 9.350 2.660 ;
        RECT  8.710 2.420 8.950 4.470 ;
        RECT  8.710 4.230 11.510 4.470 ;
        RECT  10.710 1.620 12.660 1.860 ;
        RECT  12.420 1.620 12.660 2.640 ;
        RECT  12.030 2.400 12.660 2.640 ;
        RECT  10.710 1.620 10.950 2.730 ;
        RECT  10.070 2.490 10.950 2.730 ;
        RECT  12.030 2.400 12.270 3.430 ;
        RECT  12.030 3.190 12.620 3.430 ;
        RECT  7.830 0.980 11.080 1.220 ;
        RECT  11.940 0.980 13.610 1.220 ;
        RECT  10.840 1.140 12.180 1.380 ;
        RECT  7.830 0.980 8.150 1.710 ;
        RECT  7.380 1.320 8.120 1.720 ;
        RECT  7.380 1.320 7.620 4.140 ;
        RECT  7.060 3.900 7.620 4.140 ;
        RECT  12.940 1.470 13.180 3.580 ;
        RECT  15.270 2.430 15.510 3.580 ;
        RECT  12.940 3.340 15.510 3.580 ;
        RECT  13.210 3.340 13.450 4.060 ;
        RECT  12.830 3.820 13.450 4.060 ;
        RECT  15.040 1.010 16.230 1.250 ;
        RECT  13.960 1.130 15.280 1.370 ;
        RECT  15.990 1.010 16.230 1.710 ;
        RECT  15.990 1.470 17.340 1.710 ;
        RECT  13.960 1.130 14.200 1.810 ;
        RECT  13.420 1.570 14.200 1.810 ;
        RECT  13.420 1.570 13.660 3.100 ;
        RECT  13.420 2.860 14.010 3.100 ;
        RECT  14.720 1.630 15.730 1.870 ;
        RECT  15.490 1.630 15.730 2.190 ;
        RECT  15.490 1.950 17.540 2.190 ;
        RECT  14.720 1.630 14.960 2.350 ;
        RECT  14.070 2.110 14.960 2.350 ;
        RECT  17.300 2.040 19.810 2.460 ;
        RECT  15.790 1.950 16.030 3.610 ;
    END
END decfq4

MACRO decfq2
    CLASS CORE ;
    FOREIGN decfq2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.490 2.580 14.730 3.410 ;
        RECT  14.060 2.580 14.730 3.020 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.191  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.220 5.660 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.086  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.040 3.700 3.860 3.990 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.232  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.700 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.334  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.660 2.020 16.180 2.460 ;
        RECT  15.660 1.470 15.900 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.800 5.600 ;
        RECT  16.330 4.130 16.570 5.600 ;
        RECT  15.000 4.130 15.240 5.600 ;
        RECT  13.350 4.710 13.750 5.600 ;
        RECT  9.490 4.340 10.430 5.600 ;
        RECT  5.820 4.400 6.060 5.600 ;
        RECT  4.600 4.400 4.840 5.600 ;
        RECT  1.690 4.710 2.170 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.800 0.740 ;
        RECT  16.330 0.000 16.570 1.300 ;
        RECT  14.990 0.000 15.230 1.300 ;
        RECT  12.540 0.000 12.930 0.890 ;
        RECT  9.950 0.000 10.190 1.760 ;
        RECT  5.900 0.000 6.300 0.890 ;
        RECT  4.430 0.000 4.830 0.890 ;
        RECT  1.620 0.000 2.020 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 2.450 1.650 2.690 ;
        RECT  0.820 1.710 1.060 3.450 ;
        RECT  2.440 1.470 2.680 3.450 ;
        RECT  0.850 1.060 1.430 1.370 ;
        RECT  0.850 1.130 2.130 1.370 ;
        RECT  1.890 1.130 2.130 3.460 ;
        RECT  1.550 3.220 2.130 3.460 ;
        RECT  1.550 3.220 1.790 4.470 ;
        RECT  0.920 4.230 2.650 4.470 ;
        RECT  2.410 4.380 3.250 4.620 ;
        RECT  3.920 1.610 4.160 3.460 ;
        RECT  5.130 1.640 6.250 1.880 ;
        RECT  6.010 2.570 6.460 2.970 ;
        RECT  6.010 1.640 6.250 3.500 ;
        RECT  5.130 3.260 6.250 3.500 ;
        RECT  6.490 1.610 7.020 1.930 ;
        RECT  6.780 2.140 7.140 2.540 ;
        RECT  6.490 3.270 7.020 3.670 ;
        RECT  6.780 1.610 7.020 4.120 ;
        RECT  6.780 3.880 7.340 4.120 ;
        RECT  3.180 1.130 7.510 1.370 ;
        RECT  7.270 1.130 7.510 1.930 ;
        RECT  7.380 1.720 7.620 3.000 ;
        RECT  3.180 1.130 3.420 3.450 ;
        RECT  7.270 2.760 7.510 3.620 ;
        RECT  8.750 1.470 8.990 3.620 ;
        RECT  8.670 3.300 10.430 3.620 ;
        RECT  8.010 0.990 9.690 1.230 ;
        RECT  9.450 0.990 9.690 2.380 ;
        RECT  9.450 2.140 10.680 2.380 ;
        RECT  8.010 0.990 8.250 3.620 ;
        RECT  10.610 1.550 11.160 1.790 ;
        RECT  9.620 2.670 11.160 2.910 ;
        RECT  10.920 1.550 11.160 3.640 ;
        RECT  10.910 2.670 11.160 3.640 ;
        RECT  12.130 1.610 12.690 1.850 ;
        RECT  12.130 1.610 12.370 3.330 ;
        RECT  12.130 3.090 12.630 3.330 ;
        RECT  4.410 2.520 4.650 4.160 ;
        RECT  7.640 3.860 10.710 4.100 ;
        RECT  12.390 3.090 12.630 4.120 ;
        RECT  10.530 3.880 12.630 4.120 ;
        RECT  4.410 3.920 6.540 4.160 ;
        RECT  6.300 3.920 6.540 4.600 ;
        RECT  7.640 3.860 7.880 4.600 ;
        RECT  6.300 4.360 7.880 4.600 ;
        RECT  12.610 2.090 12.850 2.800 ;
        RECT  12.610 2.560 13.110 2.800 ;
        RECT  12.870 2.560 13.110 4.600 ;
        RECT  11.380 4.360 13.110 4.600 ;
        RECT  11.430 1.130 13.390 1.370 ;
        RECT  13.150 1.130 13.390 2.320 ;
        RECT  11.430 1.130 11.670 2.100 ;
        RECT  13.150 2.080 14.340 2.320 ;
        RECT  11.650 1.860 11.890 3.640 ;
        RECT  13.710 1.540 15.420 1.780 ;
        RECT  13.350 2.710 13.590 3.890 ;
        RECT  15.180 1.540 15.420 3.890 ;
        RECT  13.350 3.650 15.420 3.890 ;
    END
END decfq2

MACRO decfq1
    CLASS CORE ;
    FOREIGN decfq1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CDN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.355  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.470 2.580 14.740 3.420 ;
        RECT  14.060 2.580 14.740 3.020 ;
        END
    END CDN
    PIN CPN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAGATEAREA 0.191  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.220 5.660 3.020 ;
        END
    END CPN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.086  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  2.040 3.700 3.860 3.990 ;
        END
    END D
    PIN ENN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.232  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.700 ;
        END
    END ENN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.265  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 2.020 16.120 2.460 ;
        RECT  15.740 1.470 16.010 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 16.240 5.600 ;
        RECT  14.990 4.140 15.230 5.600 ;
        RECT  13.370 4.710 13.770 5.600 ;
        RECT  9.490 4.340 10.430 5.600 ;
        RECT  5.820 4.400 6.060 5.600 ;
        RECT  4.600 4.400 4.840 5.600 ;
        RECT  1.690 4.710 2.170 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 16.240 0.740 ;
        RECT  14.990 0.000 15.230 1.300 ;
        RECT  12.540 0.000 12.930 0.890 ;
        RECT  9.950 0.000 10.190 1.760 ;
        RECT  5.900 0.000 6.300 0.890 ;
        RECT  4.430 0.000 4.830 0.890 ;
        RECT  1.620 0.000 2.020 0.890 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.820 2.450 1.650 2.690 ;
        RECT  0.820 1.710 1.060 3.450 ;
        RECT  2.440 1.470 2.680 3.450 ;
        RECT  0.850 1.060 1.430 1.370 ;
        RECT  0.850 1.130 2.130 1.370 ;
        RECT  1.890 1.130 2.130 3.460 ;
        RECT  1.550 3.220 2.130 3.460 ;
        RECT  1.550 3.220 1.790 4.470 ;
        RECT  0.920 4.230 2.650 4.470 ;
        RECT  2.410 4.380 3.250 4.620 ;
        RECT  3.920 1.610 4.160 3.460 ;
        RECT  5.130 1.640 6.250 1.880 ;
        RECT  6.010 2.570 6.460 2.970 ;
        RECT  6.010 1.640 6.250 3.500 ;
        RECT  5.130 3.260 6.250 3.500 ;
        RECT  6.490 1.610 7.020 1.930 ;
        RECT  6.780 2.140 7.140 2.540 ;
        RECT  6.490 3.270 7.020 3.670 ;
        RECT  6.780 1.610 7.020 4.120 ;
        RECT  6.780 3.880 7.340 4.120 ;
        RECT  3.180 1.130 7.510 1.370 ;
        RECT  7.270 1.130 7.510 1.930 ;
        RECT  7.380 1.720 7.620 3.000 ;
        RECT  3.180 1.130 3.420 3.450 ;
        RECT  7.270 2.760 7.510 3.620 ;
        RECT  8.750 1.470 8.990 3.620 ;
        RECT  8.670 3.300 10.430 3.620 ;
        RECT  8.010 0.990 9.690 1.230 ;
        RECT  9.450 0.990 9.690 2.380 ;
        RECT  9.450 2.140 10.680 2.380 ;
        RECT  8.010 0.990 8.250 3.620 ;
        RECT  10.610 1.550 11.160 1.790 ;
        RECT  9.620 2.670 11.160 2.910 ;
        RECT  10.920 1.550 11.160 3.640 ;
        RECT  10.910 2.670 11.160 3.640 ;
        RECT  12.130 1.610 12.690 1.850 ;
        RECT  12.130 1.610 12.370 3.330 ;
        RECT  12.130 3.090 12.630 3.330 ;
        RECT  4.410 2.520 4.650 4.160 ;
        RECT  7.640 3.860 10.710 4.100 ;
        RECT  12.390 3.090 12.630 4.120 ;
        RECT  10.530 3.880 12.630 4.120 ;
        RECT  4.410 3.920 6.540 4.160 ;
        RECT  6.300 3.920 6.540 4.600 ;
        RECT  7.640 3.860 7.880 4.600 ;
        RECT  6.300 4.360 7.880 4.600 ;
        RECT  12.610 2.090 12.850 2.800 ;
        RECT  12.610 2.560 13.110 2.800 ;
        RECT  12.870 2.560 13.110 4.600 ;
        RECT  11.380 4.360 13.110 4.600 ;
        RECT  11.430 1.130 13.390 1.370 ;
        RECT  13.150 1.130 13.390 2.320 ;
        RECT  11.430 1.130 11.670 2.100 ;
        RECT  13.150 2.080 14.340 2.320 ;
        RECT  11.650 1.860 11.890 3.640 ;
        RECT  13.710 1.540 15.500 1.780 ;
        RECT  13.350 2.710 13.590 3.900 ;
        RECT  15.260 1.540 15.500 3.900 ;
        RECT  13.350 3.660 15.500 3.900 ;
    END
END decfq1

MACRO cload1
    CLASS CORE ;
    FOREIGN cload1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.020 0.720 2.490 ;
        END
    END I
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 1.680 5.600 ;
        RECT  0.140 4.180 1.290 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 1.680 0.740 ;
        RECT  0.150 0.000 1.290 1.420 ;
        END
    END VSS
END cload1

MACRO clk2d2
    CLASS CORE ;
    FOREIGN clk2d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN C
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.366  LAYER M1  ;
        ANTENNAGATEAREA 0.250  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.740 2.580 11.160 2.820 ;
        RECT  9.740 2.580 10.580 3.020 ;
        RECT  10.270 1.420 10.510 3.020 ;
        RECT  9.790 1.420 10.510 1.660 ;
        RECT  9.740 2.580 9.980 3.520 ;
        END
    END C
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.344  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 1.860 5.540 2.260 ;
        RECT  4.540 1.860 4.980 2.460 ;
        RECT  4.430 2.980 4.830 3.380 ;
        RECT  4.540 1.860 4.830 3.380 ;
        END
    END CLK
    PIN CN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.358  LAYER M1  ;
        ANTENNAGATEAREA 0.189  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.790 1.670 2.070 1.910 ;
        RECT  0.790 3.200 1.890 3.440 ;
        RECT  0.790 1.670 1.060 3.440 ;
        RECT  0.640 2.260 1.060 3.020 ;
        END
    END CN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.760 5.600 ;
        RECT  10.480 4.340 10.720 5.600 ;
        RECT  9.000 4.340 9.240 5.600 ;
        RECT  6.760 3.750 7.000 5.600 ;
        RECT  5.950 4.780 6.420 5.600 ;
        RECT  4.260 4.200 4.500 5.600 ;
        RECT  2.050 4.530 2.450 5.600 ;
        RECT  0.540 4.590 0.940 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.760 0.740 ;
        RECT  10.560 0.000 10.960 1.010 ;
        RECT  8.990 0.000 9.230 1.350 ;
        RECT  6.510 0.000 6.750 1.420 ;
        RECT  4.890 0.000 5.130 1.140 ;
        RECT  2.330 0.000 2.570 1.330 ;
        RECT  0.980 0.000 1.220 1.190 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.000 0.550 1.930 ;
        RECT  0.150 1.000 0.400 3.670 ;
        RECT  0.150 3.350 0.550 3.670 ;
        RECT  2.810 1.010 3.450 1.250 ;
        RECT  2.810 1.010 3.050 2.440 ;
        RECT  1.960 2.200 3.050 2.440 ;
        RECT  2.610 2.200 2.850 3.620 ;
        RECT  2.610 3.380 3.230 3.620 ;
        RECT  3.340 1.660 3.580 3.160 ;
        RECT  3.470 2.920 3.710 4.540 ;
        RECT  3.470 4.140 3.840 4.540 ;
        RECT  2.690 4.220 3.840 4.540 ;
        RECT  5.660 1.000 5.900 1.620 ;
        RECT  3.950 1.380 5.900 1.620 ;
        RECT  3.830 2.190 4.230 2.590 ;
        RECT  5.190 2.790 6.490 3.030 ;
        RECT  3.950 1.380 4.190 3.860 ;
        RECT  3.950 3.620 5.430 3.860 ;
        RECT  5.190 2.790 5.430 4.020 ;
        RECT  4.920 3.620 5.430 4.020 ;
        RECT  6.050 1.990 6.970 2.230 ;
        RECT  6.730 2.610 7.570 2.850 ;
        RECT  6.730 1.990 6.970 3.510 ;
        RECT  6.020 3.270 6.970 3.510 ;
        RECT  6.020 3.270 6.260 3.820 ;
        RECT  7.810 1.020 8.310 1.340 ;
        RECT  7.810 1.020 8.050 3.530 ;
        RECT  7.500 3.290 8.050 3.530 ;
        RECT  7.500 3.290 7.740 4.540 ;
        RECT  7.500 4.300 8.760 4.540 ;
        RECT  8.290 1.750 8.760 2.210 ;
        RECT  8.290 1.970 9.950 2.210 ;
        RECT  8.290 1.750 8.640 3.520 ;
        RECT  11.210 1.750 11.640 2.080 ;
        RECT  11.400 1.750 11.640 3.520 ;
        RECT  11.080 3.120 11.640 3.520 ;
        RECT  11.080 3.120 11.380 4.540 ;
    END
END clk2d2

MACRO cg01d4
    CLASS CORE ;
    FOREIGN cg01d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.440 3.650 2.840 ;
        RECT  2.860 2.020 3.320 2.840 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.907  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.940 2.440 4.980 2.840 ;
        RECT  4.540 2.020 4.980 2.840 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.220 2.080 6.600 3.020 ;
        RECT  6.140 2.080 6.600 2.480 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.060  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.010 4.360 2.590 4.600 ;
        RECT  0.330 1.360 2.260 1.800 ;
        RECT  2.010 3.600 2.250 4.600 ;
        RECT  0.780 3.600 2.250 4.000 ;
        RECT  0.780 1.360 1.180 4.000 ;
        RECT  0.470 1.360 1.180 2.460 ;
        END
    END CO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  4.230 4.460 4.630 5.600 ;
        RECT  2.830 3.560 3.070 5.600 ;
        RECT  1.530 4.620 1.770 5.600 ;
        RECT  0.230 3.050 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  4.230 0.000 4.630 0.890 ;
        RECT  2.830 0.000 3.070 1.580 ;
        RECT  1.110 0.000 1.510 1.120 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.420 2.060 2.620 2.500 ;
        RECT  2.380 2.060 2.620 3.320 ;
        RECT  5.510 1.460 5.750 3.510 ;
        RECT  2.380 3.080 3.710 3.320 ;
        RECT  3.460 3.190 5.830 3.430 ;
        RECT  5.510 3.190 5.830 3.510 ;
        RECT  3.580 1.130 6.490 1.220 ;
        RECT  4.880 0.980 6.490 1.220 ;
        RECT  3.570 1.170 5.120 1.370 ;
        RECT  6.250 0.980 6.490 1.720 ;
        RECT  3.570 1.170 3.810 1.780 ;
        RECT  3.490 3.810 6.570 4.050 ;
    END
END cg01d4

MACRO cg01d2
    CLASS CORE ;
    FOREIGN cg01d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.020 0.800 2.460 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 1.820 2.460 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.331  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.160 2.020 2.780 2.460 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.162  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.350 3.130 5.460 3.370 ;
        RECT  5.100 1.850 5.460 3.370 ;
        RECT  4.350 1.850 5.460 2.090 ;
        END
    END CO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  5.000 4.130 5.240 5.600 ;
        RECT  3.690 3.730 3.930 5.600 ;
        RECT  0.970 3.730 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  5.090 0.000 5.330 1.590 ;
        RECT  3.690 0.000 3.930 1.590 ;
        RECT  0.900 0.000 1.300 1.030 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.130 2.070 3.370 ;
        RECT  0.150 1.410 2.070 1.650 ;
        RECT  2.410 1.540 3.260 1.780 ;
        RECT  3.020 2.380 4.420 2.620 ;
        RECT  3.020 1.540 3.260 3.370 ;
        RECT  2.410 3.130 3.260 3.370 ;
    END
END cg01d2

MACRO cg01d1
    CLASS CORE ;
    FOREIGN cg01d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.140 0.800 2.590 ;
        RECT  0.120 2.140 0.500 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 1.820 2.520 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.160 2.020 2.660 2.520 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.220  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 3.100 4.750 3.500 ;
        RECT  4.510 1.770 4.750 3.500 ;
        RECT  4.350 1.770 4.750 2.090 ;
        END
    END CO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.690 3.760 3.930 5.600 ;
        RECT  0.970 3.740 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.690 0.000 3.930 1.860 ;
        RECT  0.980 0.000 1.220 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.260 2.070 3.500 ;
        RECT  0.150 1.540 2.070 1.780 ;
        RECT  2.410 1.540 3.140 1.780 ;
        RECT  2.900 2.600 4.260 2.840 ;
        RECT  2.900 1.540 3.140 3.370 ;
        RECT  2.410 3.130 3.140 3.370 ;
    END
END cg01d1

MACRO cg01d0
    CLASS CORE ;
    FOREIGN cg01d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.250 1.010 2.490 ;
        RECT  0.140 2.020 0.420 2.490 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.100 1.780 2.570 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.120 2.020 2.770 2.570 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.632  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.430 2.700 4.900 3.450 ;
        RECT  4.440 1.580 4.900 3.450 ;
        RECT  4.430 1.580 4.900 1.980 ;
        END
    END CO
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.690 3.380 3.930 5.600 ;
        RECT  0.970 3.830 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.690 0.000 3.930 1.860 ;
        RECT  0.980 0.000 1.220 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.160 2.030 3.400 ;
        RECT  0.150 1.540 2.070 1.780 ;
        RECT  2.410 1.540 3.250 1.780 ;
        RECT  3.010 2.340 4.200 2.580 ;
        RECT  3.010 1.540 3.250 3.370 ;
        RECT  2.370 3.130 3.250 3.370 ;
    END
END cg01d0

MACRO buftda
    CLASS CORE ;
    FOREIGN buftda 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.401  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.410 2.210 1.060 3.020 ;
        END
    END EN
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.553  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  3.090 2.770 3.500 3.220 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.290 3.740 8.590 4.390 ;
        RECT  7.810 1.210 8.590 4.390 ;
        RECT  4.270 1.210 8.590 1.710 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.450 4.620 7.850 5.600 ;
        RECT  6.150 4.620 6.550 5.600 ;
        RECT  4.850 4.620 5.250 5.600 ;
        RECT  3.540 4.620 3.940 5.600 ;
        RECT  0.980 3.940 1.220 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.430 0.000 7.830 0.980 ;
        RECT  6.130 0.000 6.530 0.980 ;
        RECT  4.830 0.000 5.230 0.980 ;
        RECT  3.530 0.000 3.930 0.980 ;
        RECT  0.970 0.000 1.210 1.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.190 0.470 1.970 ;
        RECT  0.230 1.730 1.540 1.970 ;
        RECT  1.300 1.730 1.540 3.500 ;
        RECT  0.240 3.260 1.540 3.500 ;
        RECT  0.240 3.260 0.480 4.210 ;
        RECT  1.630 1.100 3.330 1.430 ;
        RECT  2.910 1.100 3.330 2.340 ;
        RECT  2.910 1.940 5.380 2.340 ;
        RECT  2.330 2.290 3.190 2.540 ;
        RECT  4.090 1.940 5.380 2.550 ;
        RECT  2.330 2.290 2.730 3.810 ;
        RECT  1.780 1.660 2.630 2.060 ;
        RECT  5.850 2.590 7.200 3.170 ;
        RECT  4.090 2.780 5.920 3.180 ;
        RECT  4.090 2.780 4.490 3.500 ;
        RECT  3.740 3.260 4.490 3.500 ;
        RECT  3.740 3.260 4.060 3.990 ;
        RECT  2.960 3.590 4.060 3.990 ;
        RECT  1.780 1.660 2.100 4.410 ;
        RECT  1.640 3.990 2.100 4.410 ;
        RECT  2.960 3.590 3.360 4.410 ;
        RECT  1.640 4.040 3.360 4.410 ;
    END
END buftda

MACRO buftd7
    CLASS CORE ;
    FOREIGN buftd7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.401  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.410 2.210 1.060 3.020 ;
        END
    END EN
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.554  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  3.090 2.770 3.500 3.220 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.626  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.890 3.740 7.290 4.060 ;
        RECT  6.970 3.660 7.290 4.060 ;
        RECT  6.860 1.370 7.270 1.770 ;
        RECT  6.970 1.370 7.210 4.060 ;
        RECT  6.220 1.440 7.210 1.900 ;
        RECT  4.290 3.740 7.290 3.980 ;
        RECT  4.270 1.440 7.270 1.680 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  6.150 4.620 6.550 5.600 ;
        RECT  4.850 4.620 5.250 5.600 ;
        RECT  3.540 4.620 3.940 5.600 ;
        RECT  0.980 3.940 1.220 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.130 0.000 6.530 0.980 ;
        RECT  4.830 0.000 5.230 0.980 ;
        RECT  3.520 0.000 3.920 0.980 ;
        RECT  0.970 0.000 1.210 1.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.190 0.470 1.970 ;
        RECT  0.230 1.730 1.540 1.970 ;
        RECT  1.300 1.730 1.540 3.500 ;
        RECT  0.240 3.260 1.540 3.500 ;
        RECT  0.240 3.260 0.480 4.210 ;
        RECT  1.630 1.170 3.330 1.410 ;
        RECT  2.910 1.170 3.330 2.340 ;
        RECT  2.910 2.100 4.420 2.340 ;
        RECT  2.330 2.290 3.150 2.530 ;
        RECT  2.330 2.290 2.570 3.810 ;
        RECT  1.780 1.810 2.630 2.050 ;
        RECT  4.800 2.590 5.040 3.500 ;
        RECT  3.740 3.260 5.040 3.500 ;
        RECT  3.740 3.260 3.980 3.830 ;
        RECT  2.950 3.590 3.980 3.830 ;
        RECT  1.780 1.810 2.020 4.410 ;
        RECT  1.640 3.990 2.020 4.410 ;
        RECT  2.950 3.590 3.350 4.410 ;
        RECT  1.640 4.090 3.350 4.410 ;
    END
END buftd7

MACRO buftd4
    CLASS CORE ;
    FOREIGN buftd4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.401  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.410 2.210 1.060 3.020 ;
        END
    END EN
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.506  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  3.090 2.770 3.500 3.220 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.140  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.290 3.740 6.010 3.980 ;
        RECT  5.690 1.440 6.010 3.980 ;
        RECT  5.100 1.440 6.010 1.900 ;
        RECT  4.310 1.440 6.010 1.680 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.850 4.620 5.250 5.600 ;
        RECT  3.540 4.620 3.940 5.600 ;
        RECT  0.980 3.940 1.220 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.870 0.000 5.270 0.980 ;
        RECT  3.570 0.000 3.970 0.980 ;
        RECT  0.970 0.000 1.210 1.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.190 0.470 1.970 ;
        RECT  0.230 1.730 1.540 1.970 ;
        RECT  1.300 1.730 1.540 3.500 ;
        RECT  0.240 3.260 1.540 3.500 ;
        RECT  0.240 3.260 0.480 4.210 ;
        RECT  1.630 1.170 3.330 1.410 ;
        RECT  2.910 1.170 3.330 2.340 ;
        RECT  2.910 2.100 4.460 2.340 ;
        RECT  2.330 2.290 3.150 2.530 ;
        RECT  2.330 2.290 2.570 3.810 ;
        RECT  1.780 1.810 2.630 2.050 ;
        RECT  4.800 2.590 5.040 3.500 ;
        RECT  3.740 3.260 5.040 3.500 ;
        RECT  3.740 3.260 3.980 3.830 ;
        RECT  2.950 3.590 3.980 3.830 ;
        RECT  1.780 1.810 2.020 4.440 ;
        RECT  1.640 3.990 2.020 4.440 ;
        RECT  2.950 3.590 3.350 4.330 ;
        RECT  1.640 4.090 3.350 4.330 ;
        RECT  1.640 4.090 2.040 4.440 ;
    END
END buftd4

MACRO buftd2
    CLASS CORE ;
    FOREIGN buftd2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.410 2.210 1.060 3.020 ;
        END
    END EN
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.508  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  3.330 2.920 3.730 3.350 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.259  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.450 3.810 5.460 4.050 ;
        RECT  5.180 1.300 5.460 4.050 ;
        RECT  5.100 1.300 5.460 1.900 ;
        RECT  4.410 1.300 5.460 1.540 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  5.040 4.620 5.440 5.600 ;
        RECT  3.670 4.620 4.070 5.600 ;
        RECT  0.980 3.940 1.220 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  5.010 0.000 5.410 0.980 ;
        RECT  3.670 0.000 4.070 0.980 ;
        RECT  0.970 0.000 1.210 1.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.190 0.470 1.970 ;
        RECT  0.230 1.730 1.710 1.970 ;
        RECT  1.470 1.730 1.710 3.500 ;
        RECT  0.240 3.260 1.710 3.500 ;
        RECT  0.240 3.260 0.480 4.110 ;
        RECT  1.980 1.810 2.670 2.050 ;
        RECT  4.100 2.950 4.340 3.590 ;
        RECT  1.980 1.810 2.220 4.230 ;
        RECT  3.970 3.350 4.210 4.060 ;
        RECT  3.080 3.820 4.210 4.060 ;
        RECT  1.640 3.990 3.480 4.230 ;
        RECT  1.670 1.170 3.420 1.410 ;
        RECT  2.910 1.170 3.420 2.070 ;
        RECT  2.910 1.830 4.560 2.070 ;
        RECT  2.910 1.170 3.150 2.530 ;
        RECT  2.460 2.290 3.150 2.530 ;
        RECT  2.460 2.290 2.700 3.710 ;
    END
END buftd2

MACRO buftd1
    CLASS CORE ;
    FOREIGN buftd1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.401  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.540 1.060 3.020 ;
        END
    END EN
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.320 2.860 3.860 3.580 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.490 4.280 4.920 4.600 ;
        RECT  4.680 1.000 4.920 4.600 ;
        RECT  4.400 1.000 4.920 1.900 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.740 4.480 3.980 5.600 ;
        RECT  0.970 3.960 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.660 0.000 4.060 1.070 ;
        RECT  0.970 0.000 1.210 1.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.190 0.470 1.970 ;
        RECT  0.230 1.730 1.700 1.970 ;
        RECT  1.460 1.730 1.700 3.610 ;
        RECT  0.230 3.370 1.700 3.610 ;
        RECT  0.230 3.370 0.470 4.130 ;
        RECT  1.970 1.810 2.630 2.050 ;
        RECT  1.970 1.810 2.210 4.220 ;
        RECT  3.070 3.820 4.340 4.060 ;
        RECT  4.100 2.860 4.340 4.060 ;
        RECT  1.630 3.980 3.470 4.220 ;
        RECT  1.630 1.170 3.390 1.410 ;
        RECT  3.070 2.140 4.400 2.380 ;
        RECT  3.070 1.170 3.390 2.530 ;
        RECT  2.450 2.290 3.390 2.530 ;
        RECT  2.450 2.290 2.690 3.740 ;
    END
END buftd1

MACRO buffda
    CLASS CORE ;
    FOREIGN buffda 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.178  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.300 1.080 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.095  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.790 3.130 7.160 3.630 ;
        RECT  4.190 1.770 7.160 3.630 ;
        RECT  3.030 1.770 7.160 2.270 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  5.980 4.620 6.380 5.600 ;
        RECT  4.650 4.620 5.050 5.600 ;
        RECT  3.350 4.620 3.750 5.600 ;
        RECT  2.050 4.620 2.450 5.600 ;
        RECT  0.800 3.870 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.730 0.000 7.130 0.980 ;
        RECT  5.250 0.000 5.650 0.980 ;
        RECT  3.770 0.000 4.170 0.980 ;
        RECT  2.290 0.000 2.690 0.970 ;
        RECT  0.920 0.000 1.320 1.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.650 2.090 2.050 ;
        RECT  1.690 2.500 3.960 2.900 ;
        RECT  1.690 1.650 2.090 3.640 ;
        RECT  0.150 3.250 2.090 3.640 ;
    END
END buffda

MACRO buffd7
    CLASS CORE ;
    FOREIGN buffd7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.780  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.520 2.020 1.060 2.700 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.351  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.940 3.050 5.350 3.450 ;
        RECT  4.540 2.580 4.980 3.400 ;
        RECT  4.540 1.460 4.780 3.400 ;
        RECT  2.230 3.160 5.350 3.400 ;
        RECT  2.230 1.460 4.780 1.700 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.240 4.610 4.640 5.600 ;
        RECT  2.820 4.610 3.220 5.600 ;
        RECT  1.520 4.560 1.920 5.600 ;
        RECT  0.280 3.860 0.520 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.450 0.000 4.850 0.980 ;
        RECT  2.970 0.000 3.370 0.980 ;
        RECT  1.490 0.000 1.890 0.970 ;
        RECT  0.230 0.000 0.470 1.710 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.890 1.540 1.540 1.780 ;
        RECT  1.300 2.600 2.260 2.840 ;
        RECT  1.300 1.540 1.540 3.370 ;
        RECT  0.770 3.130 1.540 3.370 ;
    END
END buffd7

MACRO buffd4
    CLASS CORE ;
    FOREIGN buffd4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.582  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.470 2.370 1.060 2.830 ;
        RECT  0.620 2.020 1.060 2.830 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.410 2.560 3.910 2.800 ;
        RECT  3.670 0.980 3.910 2.800 ;
        RECT  2.030 1.270 3.910 1.510 ;
        RECT  3.510 0.980 3.910 1.510 ;
        RECT  3.410 2.560 3.650 4.280 ;
        RECT  2.020 3.070 3.650 3.470 ;
        RECT  2.300 3.070 2.740 4.140 ;
        RECT  2.030 0.980 2.430 1.510 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.920 3.050 4.320 5.600 ;
        RECT  2.760 4.620 3.160 5.600 ;
        RECT  1.460 4.490 1.860 5.600 ;
        RECT  0.150 3.750 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  2.770 0.000 3.170 0.980 ;
        RECT  1.290 0.000 1.690 1.150 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.540 1.780 ;
        RECT  1.300 1.750 3.250 2.150 ;
        RECT  1.300 1.540 1.540 3.390 ;
        RECT  0.720 3.150 1.540 3.390 ;
    END
END buffd4

MACRO buffd3
    CLASS CORE ;
    FOREIGN buffd3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.300 0.540 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.571  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.550 2.120 3.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  2.240 4.620 2.640 5.600 ;
        RECT  1.000 4.200 1.240 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  2.320 0.000 2.560 1.180 ;
        RECT  1.020 0.000 1.260 1.390 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.660 1.320 1.900 ;
        RECT  1.080 2.300 1.520 2.700 ;
        RECT  1.080 1.660 1.320 3.950 ;
        RECT  0.150 3.710 1.320 3.950 ;
    END
END buffd3

MACRO buffd2
    CLASS CORE ;
    FOREIGN buffd2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.850 1.060 2.460 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.550  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.020 2.680 2.460 ;
        RECT  1.680 3.250 2.590 3.490 ;
        RECT  2.300 1.580 2.590 3.490 ;
        RECT  1.710 1.580 2.590 1.820 ;
        RECT  1.710 1.090 1.950 1.820 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.330 4.110 2.570 5.600 ;
        RECT  0.800 3.730 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.450 0.000 2.690 1.320 ;
        RECT  0.970 0.000 1.210 1.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.210 0.550 1.610 ;
        RECT  1.500 2.060 1.900 2.940 ;
        RECT  1.200 2.700 1.900 2.940 ;
        RECT  0.120 1.210 0.360 3.450 ;
        RECT  1.200 2.700 1.440 3.370 ;
        RECT  0.120 3.130 1.440 3.370 ;
        RECT  0.120 3.050 0.490 3.450 ;
    END
END buffd2

MACRO buffd1
    CLASS CORE ;
    FOREIGN buffd1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.020 0.540 2.590 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.014  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.550 2.120 3.580 ;
        RECT  1.750 1.550 2.120 1.950 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.240 5.600 ;
        RECT  1.170 4.050 1.410 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.240 0.740 ;
        RECT  1.140 0.000 1.380 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.270 1.540 1.320 1.780 ;
        RECT  1.080 2.080 1.520 2.480 ;
        RECT  1.080 1.540 1.320 3.370 ;
        RECT  0.270 3.130 1.320 3.370 ;
    END
END buffd1

MACRO bufbdk
    CLASS CORE ;
    FOREIGN bufbdk 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.177  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.360 2.400 1.280 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 13.276  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.330 1.220 12.820 3.580 ;
        RECT  2.750 2.510 12.820 3.550 ;
        RECT  4.120 1.220 12.820 3.550 ;
        RECT  3.110 1.220 12.820 1.650 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 13.440 5.600 ;
        RECT  12.650 4.620 13.050 5.600 ;
        RECT  11.300 4.590 11.700 5.600 ;
        RECT  10.000 4.580 10.400 5.600 ;
        RECT  8.700 4.600 9.100 5.600 ;
        RECT  7.400 4.590 7.800 5.600 ;
        RECT  6.100 4.590 6.500 5.600 ;
        RECT  4.800 4.590 5.200 5.600 ;
        RECT  3.500 4.600 3.900 5.600 ;
        RECT  2.050 4.580 2.450 5.600 ;
        RECT  0.720 4.160 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 13.440 0.740 ;
        RECT  12.750 0.000 13.150 0.980 ;
        RECT  11.270 0.000 11.670 0.980 ;
        RECT  9.770 0.000 10.170 0.980 ;
        RECT  8.290 0.000 8.690 0.980 ;
        RECT  6.810 0.000 7.210 0.980 ;
        RECT  5.330 0.000 5.730 0.980 ;
        RECT  3.850 0.000 4.250 0.980 ;
        RECT  2.370 0.000 2.770 1.480 ;
        RECT  0.890 0.000 1.290 1.520 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.140 1.090 0.550 2.170 ;
        RECT  0.140 1.770 2.030 2.170 ;
        RECT  1.630 1.090 2.030 2.170 ;
        RECT  1.670 1.880 3.890 2.280 ;
        RECT  1.670 1.880 2.070 3.790 ;
        RECT  0.140 3.390 2.070 3.790 ;
    END
END bufbdk

MACRO bufbdf
    CLASS CORE ;
    FOREIGN bufbdf 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.871  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.910 2.580 1.620 3.020 ;
        RECT  0.910 2.040 1.310 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 10.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.760 2.630 10.240 4.060 ;
        RECT  4.120 1.240 10.240 4.060 ;
        RECT  3.110 1.240 10.240 1.770 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  10.000 4.600 10.400 5.600 ;
        RECT  8.700 4.600 9.100 5.600 ;
        RECT  7.400 4.600 7.800 5.600 ;
        RECT  6.100 4.600 6.500 5.600 ;
        RECT  4.800 4.600 5.200 5.600 ;
        RECT  3.500 4.600 3.900 5.600 ;
        RECT  2.150 4.600 2.550 5.600 ;
        RECT  0.800 4.080 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  9.890 0.000 10.290 0.980 ;
        RECT  8.290 0.000 8.690 0.980 ;
        RECT  6.810 0.000 7.210 0.980 ;
        RECT  5.330 0.000 5.730 0.980 ;
        RECT  3.850 0.000 4.250 0.980 ;
        RECT  2.450 0.000 2.690 1.510 ;
        RECT  0.970 0.000 1.210 1.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.630 1.060 2.030 2.340 ;
        RECT  1.960 2.000 3.890 2.400 ;
        RECT  0.150 1.060 0.550 3.760 ;
        RECT  1.960 2.000 2.360 3.760 ;
        RECT  0.150 3.360 2.360 3.760 ;
    END
END bufbdf

MACRO bufbda
    CLASS CORE ;
    FOREIGN bufbda 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.121  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.580 1.910 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.280  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.870 3.000 8.540 3.600 ;
        RECT  4.250 1.480 6.420 3.600 ;
        RECT  4.640 1.440 5.040 3.600 ;
        RECT  3.270 1.480 6.420 2.080 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  8.880 4.560 9.280 5.600 ;
        RECT  7.550 4.560 7.950 5.600 ;
        RECT  6.250 4.560 6.650 5.600 ;
        RECT  4.950 4.560 5.350 5.600 ;
        RECT  3.690 4.380 3.930 5.600 ;
        RECT  2.390 4.180 2.630 5.600 ;
        RECT  0.820 4.180 1.060 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  6.790 0.000 7.190 0.980 ;
        RECT  5.210 0.000 5.610 0.980 ;
        RECT  3.790 0.000 4.190 0.980 ;
        RECT  2.460 0.000 2.860 0.980 ;
        RECT  1.030 0.000 1.270 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 2.550 1.940 ;
        RECT  2.150 1.540 2.550 2.760 ;
        RECT  2.150 2.360 4.020 2.760 ;
        RECT  0.150 1.540 0.550 3.650 ;
        RECT  0.150 3.250 1.850 3.650 ;
    END
END bufbda

MACRO bufbd7
    CLASS CORE ;
    FOREIGN bufbd7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.138  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.580 1.910 3.030 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.957  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.980 3.220 7.330 3.460 ;
        RECT  3.050 1.460 6.230 1.700 ;
        RECT  3.410 1.460 3.920 1.910 ;
        RECT  3.500 1.460 3.780 3.460 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  6.450 4.370 6.690 5.600 ;
        RECT  5.150 4.370 5.390 5.600 ;
        RECT  3.810 4.370 4.050 5.600 ;
        RECT  2.240 4.180 2.480 5.600 ;
        RECT  0.820 4.180 1.060 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  5.060 0.000 5.460 0.990 ;
        RECT  3.870 0.000 4.110 1.130 ;
        RECT  2.540 0.000 2.780 1.130 ;
        RECT  1.020 0.000 1.260 1.330 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.620 2.390 1.860 ;
        RECT  0.150 1.620 0.550 2.020 ;
        RECT  2.150 1.620 2.390 2.830 ;
        RECT  2.150 2.590 3.130 2.830 ;
        RECT  0.230 1.620 0.550 3.540 ;
        RECT  0.150 3.140 0.550 3.540 ;
        RECT  0.150 3.300 1.850 3.540 ;
    END
END bufbd7

MACRO bufbd4
    CLASS CORE ;
    FOREIGN bufbd4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.538  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.470 1.340 3.020 ;
        RECT  1.000 2.440 1.340 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.988  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.370 1.130 3.770 4.440 ;
        RECT  2.060 2.580 3.770 3.020 ;
        RECT  1.890 1.220 3.770 1.460 ;
        RECT  1.890 1.130 2.290 1.460 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  2.620 3.370 3.020 5.600 ;
        RECT  1.200 4.610 1.600 5.600 ;
        RECT  0.150 3.870 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  2.630 0.000 3.030 0.980 ;
        RECT  1.150 0.000 1.550 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.290 0.550 2.020 ;
        RECT  0.150 1.780 2.710 2.020 ;
        RECT  1.580 1.780 2.710 2.180 ;
        RECT  1.580 1.780 1.820 3.520 ;
        RECT  0.720 3.280 1.820 3.520 ;
    END
END bufbd4

MACRO bufbd3
    CLASS CORE ;
    FOREIGN bufbd3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.662  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.140 0.720 2.540 ;
        RECT  0.140 2.140 0.500 3.020 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.045  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.040 3.130 3.740 3.370 ;
        RECT  2.980 1.460 3.300 3.370 ;
        RECT  2.630 1.460 3.300 1.900 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  2.860 4.090 3.100 5.600 ;
        RECT  1.560 3.910 1.800 5.600 ;
        RECT  0.230 3.910 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  3.370 0.000 3.770 1.020 ;
        RECT  2.070 0.000 2.470 1.020 ;
        RECT  1.000 0.000 1.240 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.660 1.200 1.900 ;
        RECT  0.960 2.600 2.190 2.840 ;
        RECT  0.960 1.660 1.200 3.530 ;
        RECT  0.720 3.130 1.200 3.530 ;
    END
END bufbd3

MACRO bufbd2
    CLASS CORE ;
    FOREIGN bufbd2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.506  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.480 2.370 0.720 3.020 ;
        RECT  0.120 1.790 0.500 2.610 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.303  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.240 3.830 2.640 4.230 ;
        RECT  2.370 1.440 2.610 4.230 ;
        RECT  2.110 1.440 2.610 1.680 ;
        RECT  2.110 0.980 2.350 1.680 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.810 4.620 3.210 5.600 ;
        RECT  1.740 3.100 1.980 5.600 ;
        RECT  0.150 4.110 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.770 0.000 3.170 1.080 ;
        RECT  1.290 0.000 1.690 1.080 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.300 1.180 1.540 ;
        RECT  0.940 1.370 1.210 1.610 ;
        RECT  0.970 1.920 2.100 2.320 ;
        RECT  0.970 1.370 1.210 4.060 ;
    END
END bufbd2

MACRO bufbd1
    CLASS CORE ;
    FOREIGN bufbd1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.314  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.960 1.050 2.380 ;
        RECT  0.600 1.960 0.940 2.460 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.929  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.630 3.080 2.260 3.320 ;
        RECT  2.020 1.380 2.260 3.320 ;
        RECT  1.630 1.380 2.260 1.910 ;
        RECT  1.630 3.080 1.880 3.630 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  2.190 3.910 2.430 5.600 ;
        RECT  0.800 3.910 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  0.970 0.000 1.210 1.720 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.120 1.380 0.550 1.700 ;
        RECT  1.150 2.600 1.780 2.840 ;
        RECT  0.120 1.380 0.360 3.640 ;
        RECT  1.150 2.600 1.390 3.640 ;
        RECT  0.120 3.230 1.390 3.640 ;
    END
END bufbd1

MACRO bh01d1
    CLASS CORE ;
    FOREIGN bh01d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INOUT ;
        ANTENNADIFFAREA 0.429  LAYER M1  ;
        ANTENNAGATEAREA 0.207  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.760 3.860 2.750 ;
        RECT  3.150 1.760 3.390 3.620 ;
        END
    END I
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.920 4.170 4.320 5.600 ;
        RECT  0.180 3.220 0.580 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.920 0.000 4.320 1.460 ;
        RECT  0.150 0.000 0.550 2.170 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.300 1.060 3.580 1.460 ;
        RECT  0.610 2.420 2.890 2.820 ;
        RECT  2.490 1.060 2.890 4.360 ;
        RECT  2.240 3.960 3.580 4.360 ;
    END
END bh01d1

MACRO aor31d4
    CLASS CORE ;
    FOREIGN aor31d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.540 2.800 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.090 2.580 1.540 3.210 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.392  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.780 1.900 2.110 2.550 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.350 2.020 2.720 3.210 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.291  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.390 3.900 5.090 4.300 ;
        RECT  3.470 2.060 5.010 2.300 ;
        RECT  4.770 1.620 5.010 2.300 ;
        RECT  3.640 3.700 4.420 4.300 ;
        RECT  3.640 2.060 3.880 4.300 ;
        RECT  3.470 1.620 3.710 2.300 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  3.960 4.620 4.360 5.600 ;
        RECT  2.620 4.710 3.020 5.600 ;
        RECT  1.490 4.710 1.890 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  3.960 0.000 4.360 1.330 ;
        RECT  2.580 0.000 2.980 0.890 ;
        RECT  0.230 0.000 0.470 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 3.450 2.420 3.690 ;
        RECT  0.890 1.100 2.380 1.340 ;
        RECT  2.140 1.130 3.200 1.370 ;
        RECT  2.960 2.520 3.360 2.920 ;
        RECT  2.960 1.130 3.200 3.690 ;
        RECT  2.710 3.450 3.200 3.690 ;
        RECT  2.710 3.450 2.950 4.380 ;
        RECT  0.150 4.140 2.950 4.380 ;
    END
END aor31d4

MACRO aor31d2
    CLASS CORE ;
    FOREIGN aor31d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.540 2.800 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.090 2.580 1.540 3.210 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.392  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.780 1.900 2.110 2.550 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.350 2.020 2.720 3.210 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.365  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.360 3.900 3.860 4.300 ;
        RECT  3.620 2.060 3.860 4.300 ;
        RECT  3.440 1.620 3.680 2.300 ;
        RECT  3.450 3.700 3.860 4.300 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.930 4.620 4.330 5.600 ;
        RECT  2.590 4.710 2.990 5.600 ;
        RECT  1.500 4.710 1.900 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.930 0.000 4.330 1.330 ;
        RECT  2.580 0.000 2.980 0.890 ;
        RECT  0.230 0.000 0.470 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 3.450 2.420 3.690 ;
        RECT  0.890 1.100 2.380 1.340 ;
        RECT  2.140 1.130 3.200 1.370 ;
        RECT  2.960 2.600 3.360 3.000 ;
        RECT  2.960 1.130 3.200 3.690 ;
        RECT  2.700 3.450 3.200 3.690 ;
        RECT  2.700 3.450 2.940 4.380 ;
        RECT  0.150 4.140 2.940 4.380 ;
    END
END aor31d2

MACRO aor31d1
    CLASS CORE ;
    FOREIGN aor31d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.020 0.460 2.800 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.140 1.620 3.580 ;
        RECT  1.180 2.750 1.420 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.690 2.020 2.180 2.530 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.590 3.700 3.300 4.140 ;
        RECT  2.590 2.750 2.830 4.140 ;
        RECT  2.290 2.750 2.830 3.150 ;
        END
    END B3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.143  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 2.550 3.800 3.510 ;
        RECT  3.450 1.350 3.690 3.510 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  2.880 4.380 3.120 5.600 ;
        RECT  1.440 4.710 1.860 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  2.580 0.000 2.980 0.890 ;
        RECT  0.230 0.000 0.470 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.110 3.390 2.350 4.310 ;
        RECT  0.720 4.070 2.350 4.310 ;
        RECT  0.710 1.080 2.380 1.320 ;
        RECT  2.140 1.130 3.210 1.370 ;
        RECT  0.710 1.080 0.950 2.390 ;
        RECT  2.970 1.130 3.210 2.530 ;
        RECT  0.700 2.150 0.940 3.610 ;
        RECT  0.150 3.370 0.940 3.610 ;
    END
END aor31d1

MACRO aor311d4
    CLASS CORE ;
    FOREIGN aor311d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.020 0.500 2.950 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.395  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.700 1.480 3.940 ;
        RECT  1.220 2.580 1.480 3.940 ;
        RECT  0.620 3.700 1.060 4.140 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.545  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.180 2.710 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.563  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.500 2.640 2.900 3.040 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.500 2.640 2.740 3.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.545  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.340 3.140 3.860 3.580 ;
        RECT  3.340 2.580 3.580 3.580 ;
        RECT  3.180 2.580 3.580 2.980 ;
        END
    END C3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.762  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.300 3.140 6.000 3.500 ;
        RECT  5.760 1.750 6.000 3.500 ;
        RECT  4.300 1.830 6.000 2.070 ;
        RECT  5.600 1.750 6.000 2.070 ;
        RECT  5.100 3.140 5.540 3.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.940 4.450 5.180 5.600 ;
        RECT  3.640 4.450 3.880 5.600 ;
        RECT  2.200 4.520 2.440 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.980 0.000 5.220 1.440 ;
        RECT  3.460 0.000 3.860 0.910 ;
        RECT  0.970 0.000 1.370 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.720 3.920 3.190 4.160 ;
        RECT  1.720 3.920 1.960 4.420 ;
        RECT  1.380 4.180 1.780 4.580 ;
        RECT  0.740 1.240 4.070 1.480 ;
        RECT  1.740 1.160 2.140 1.560 ;
        RECT  0.150 1.490 0.980 1.730 ;
        RECT  3.820 1.240 4.060 2.620 ;
        RECT  3.820 2.380 4.990 2.620 ;
        RECT  0.740 1.240 0.980 3.460 ;
        RECT  0.150 3.220 0.980 3.460 ;
    END
END aor311d4

MACRO aor311d2
    CLASS CORE ;
    FOREIGN aor311d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.020 0.500 2.950 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 3.140 1.540 3.580 ;
        RECT  1.220 1.920 1.460 3.580 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.750 2.300 2.100 3.020 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.430 2.020 2.670 3.040 ;
        RECT  2.340 2.020 2.670 2.460 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.910 2.580 3.220 3.020 ;
        RECT  2.910 1.960 3.180 3.020 ;
        END
    END C3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.202  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.920 3.140 4.690 3.580 ;
        RECT  4.450 1.470 4.690 3.580 ;
        RECT  3.920 1.470 4.690 1.710 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.490 4.120 4.890 5.600 ;
        RECT  3.180 4.120 3.580 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.490 0.000 4.890 1.060 ;
        RECT  3.180 0.000 3.580 1.060 ;
        RECT  0.720 0.000 1.130 1.080 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.170 3.500 3.020 3.740 ;
        RECT  2.170 3.500 2.410 4.440 ;
        RECT  1.180 4.200 2.410 4.440 ;
        RECT  0.150 1.440 3.680 1.680 ;
        RECT  3.440 1.440 3.680 2.480 ;
        RECT  3.440 2.240 4.120 2.480 ;
        RECT  0.740 1.440 0.980 3.490 ;
        RECT  0.150 3.250 0.980 3.490 ;
    END
END aor311d2

MACRO aor311d1
    CLASS CORE ;
    FOREIGN aor311d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.020 0.500 2.950 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 3.140 1.540 3.580 ;
        RECT  1.220 1.920 1.460 3.580 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.750 2.300 2.100 3.020 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.430 2.020 2.670 3.040 ;
        RECT  2.340 2.020 2.670 2.460 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.910 2.580 3.220 3.020 ;
        RECT  2.910 1.960 3.180 3.020 ;
        END
    END C3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.235  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.920 3.170 4.360 4.140 ;
        RECT  4.120 1.360 4.360 4.140 ;
        RECT  3.920 1.360 4.360 1.760 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.180 4.120 3.580 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.180 0.000 3.580 1.060 ;
        RECT  0.720 0.000 1.130 1.080 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.170 3.500 3.020 3.740 ;
        RECT  2.170 3.500 2.410 4.440 ;
        RECT  1.180 4.200 2.410 4.440 ;
        RECT  0.150 1.440 3.660 1.680 ;
        RECT  3.420 1.440 3.660 2.300 ;
        RECT  3.630 2.000 3.870 2.900 ;
        RECT  0.740 1.440 0.980 3.490 ;
        RECT  0.150 3.250 0.980 3.490 ;
    END
END aor311d1

MACRO aor22d4
    CLASS CORE ;
    FOREIGN aor22d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.340 2.050 2.580 ;
        RECT  1.650 2.070 2.050 2.580 ;
        RECT  1.180 2.340 1.620 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.412  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.770 2.020 3.300 2.470 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.700 1.370 2.100 ;
        RECT  0.620 1.460 1.280 1.900 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.140 0.630 2.540 ;
        RECT  0.120 2.140 0.500 3.020 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.819  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.200 3.700 5.910 4.140 ;
        RECT  3.930 1.770 5.790 2.170 ;
        RECT  4.900 1.770 5.140 4.140 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.770 4.620 5.170 5.600 ;
        RECT  3.460 4.620 3.860 5.600 ;
        RECT  0.800 3.980 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.730 0.000 4.970 1.420 ;
        RECT  3.040 0.000 3.280 1.420 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.260 0.550 3.740 ;
        RECT  0.150 3.500 1.780 3.740 ;
        RECT  1.460 3.500 1.780 4.380 ;
        RECT  2.840 3.190 3.080 4.040 ;
        RECT  1.460 3.800 3.080 4.040 ;
        RECT  1.460 3.800 1.860 4.380 ;
        RECT  1.490 1.100 2.530 1.340 ;
        RECT  3.630 2.520 4.570 2.950 ;
        RECT  2.290 2.710 4.570 2.950 ;
        RECT  2.290 1.100 2.530 3.450 ;
        RECT  2.020 3.050 2.530 3.450 ;
    END
END aor22d4

MACRO aor22d2
    CLASS CORE ;
    FOREIGN aor22d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.340 2.050 2.580 ;
        RECT  1.650 2.070 2.050 2.580 ;
        RECT  1.180 2.340 1.620 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.780 2.020 3.300 2.470 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.700 1.370 2.100 ;
        RECT  0.620 1.460 1.280 1.900 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.140 0.630 2.540 ;
        RECT  0.120 2.140 0.500 3.020 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.230  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.920 1.540 4.360 4.240 ;
        RECT  3.770 1.540 4.360 1.940 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.490 4.620 4.890 5.600 ;
        RECT  3.170 4.650 3.570 5.600 ;
        RECT  0.800 3.980 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.570 0.000 4.810 1.420 ;
        RECT  3.040 0.000 3.280 1.420 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.260 0.550 3.740 ;
        RECT  0.150 3.500 1.780 3.740 ;
        RECT  1.460 3.500 1.780 4.380 ;
        RECT  2.840 3.190 3.080 4.040 ;
        RECT  1.460 3.800 3.080 4.040 ;
        RECT  1.460 3.800 1.860 4.380 ;
        RECT  1.490 1.060 2.530 1.300 ;
        RECT  2.290 2.710 3.610 2.950 ;
        RECT  2.290 1.060 2.530 3.450 ;
        RECT  2.020 3.050 2.530 3.450 ;
        RECT  3.370 2.710 3.610 3.560 ;
    END
END aor22d2

MACRO aor22d1
    CLASS CORE ;
    FOREIGN aor22d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.340 2.050 2.580 ;
        RECT  1.650 2.070 2.050 2.580 ;
        RECT  1.180 2.340 1.620 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.780 2.020 3.300 2.470 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.700 1.370 2.100 ;
        RECT  0.620 1.460 1.280 1.900 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.140 0.630 2.540 ;
        RECT  0.120 2.140 0.500 3.020 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.055  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.500 4.360 4.230 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.230 4.620 3.630 5.600 ;
        RECT  0.800 3.980 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.040 0.000 3.280 1.420 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.260 0.550 3.740 ;
        RECT  0.150 3.500 1.780 3.740 ;
        RECT  1.460 3.500 1.780 4.380 ;
        RECT  2.840 3.190 3.080 4.040 ;
        RECT  1.460 3.800 3.080 4.040 ;
        RECT  1.460 3.800 1.860 4.380 ;
        RECT  1.490 1.060 2.530 1.300 ;
        RECT  2.290 2.710 3.610 2.950 ;
        RECT  2.290 1.060 2.530 3.450 ;
        RECT  2.020 3.050 2.530 3.450 ;
        RECT  3.370 2.710 3.610 3.560 ;
    END
END aor22d1

MACRO aor222d4
    CLASS CORE ;
    FOREIGN aor222d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.460 1.290 2.890 ;
        RECT  0.620 1.460 1.290 1.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.429  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.140 0.630 2.540 ;
        RECT  0.120 2.140 0.500 3.020 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.020 2.520 2.680 2.920 ;
        RECT  2.290 2.020 2.680 2.920 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.920 2.020 3.350 2.420 ;
        RECT  2.920 2.020 3.300 3.020 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.300 4.420 3.020 ;
        RECT  3.840 2.300 4.420 2.700 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.551  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.660 2.580 5.540 3.020 ;
        RECT  4.660 2.520 5.060 3.020 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.235  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.980 3.140 7.690 3.580 ;
        RECT  5.870 1.460 7.690 1.700 ;
        RECT  7.090 1.460 7.330 3.580 ;
        RECT  5.980 3.140 6.380 4.620 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  6.720 4.090 7.120 5.600 ;
        RECT  5.210 4.710 5.610 5.600 ;
        RECT  4.030 4.080 4.430 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.650 0.000 7.050 1.160 ;
        RECT  5.130 0.000 5.530 1.270 ;
        RECT  3.010 0.000 3.410 1.100 ;
        RECT  0.150 0.000 0.550 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 4.120 3.130 4.360 ;
        RECT  2.160 3.260 5.170 3.500 ;
        RECT  1.530 1.340 4.110 1.750 ;
        RECT  1.530 1.510 5.630 1.750 ;
        RECT  5.390 1.510 5.630 2.340 ;
        RECT  5.390 2.100 6.820 2.340 ;
        RECT  5.880 2.100 6.820 2.700 ;
        RECT  1.530 1.340 1.770 3.370 ;
        RECT  0.720 3.130 1.770 3.370 ;
    END
END aor222d4

MACRO aor222d2
    CLASS CORE ;
    FOREIGN aor222d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.460 1.290 2.890 ;
        RECT  0.620 1.460 1.290 1.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.429  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.140 0.630 2.540 ;
        RECT  0.120 2.140 0.500 3.020 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.449  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.020 2.520 2.680 2.920 ;
        RECT  2.290 2.020 2.680 2.920 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.920 2.020 3.350 2.420 ;
        RECT  2.920 2.020 3.300 3.020 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.020 4.420 3.020 ;
        RECT  3.960 2.020 4.420 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.670 2.580 5.540 3.020 ;
        RECT  4.670 2.110 5.070 3.020 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.217  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.160 3.050 6.660 3.580 ;
        RECT  6.260 1.460 6.500 3.580 ;
        RECT  5.870 1.460 6.500 1.700 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.730 4.090 7.130 5.600 ;
        RECT  5.390 4.090 5.790 5.600 ;
        RECT  4.030 4.150 4.430 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.670 0.000 7.070 1.270 ;
        RECT  5.130 0.000 5.530 1.270 ;
        RECT  3.010 0.000 3.410 1.100 ;
        RECT  0.150 0.000 0.550 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 4.120 3.130 4.360 ;
        RECT  2.160 3.430 5.170 3.670 ;
        RECT  1.530 1.340 4.110 1.750 ;
        RECT  1.530 1.510 5.630 1.750 ;
        RECT  5.390 1.510 5.630 2.340 ;
        RECT  5.390 1.940 6.020 2.340 ;
        RECT  1.530 1.340 1.770 3.370 ;
        RECT  0.720 3.130 1.770 3.370 ;
    END
END aor222d2

MACRO aor222d1
    CLASS CORE ;
    FOREIGN aor222d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.460 1.290 2.890 ;
        RECT  0.620 1.460 1.290 1.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.429  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.140 0.630 2.540 ;
        RECT  0.120 2.140 0.500 3.020 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.449  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.020 2.520 2.680 2.920 ;
        RECT  2.290 2.020 2.680 2.920 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.920 2.020 3.350 2.420 ;
        RECT  2.920 2.020 3.300 3.020 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.020 4.420 3.020 ;
        RECT  3.960 2.020 4.420 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.880 2.020 5.540 2.460 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.029  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 3.050 6.500 3.580 ;
        RECT  6.260 1.060 6.500 3.580 ;
        RECT  5.870 1.060 6.500 1.300 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.470 4.090 5.870 5.600 ;
        RECT  4.030 4.150 4.430 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.130 0.000 5.530 1.300 ;
        RECT  3.010 0.000 3.410 1.130 ;
        RECT  0.150 0.000 0.550 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 4.120 3.130 4.360 ;
        RECT  2.160 3.430 5.170 3.670 ;
        RECT  1.530 1.370 4.110 1.780 ;
        RECT  1.530 1.540 6.020 1.780 ;
        RECT  5.780 1.540 6.020 2.420 ;
        RECT  1.530 1.370 1.770 3.370 ;
        RECT  0.720 3.130 1.770 3.370 ;
    END
END aor222d1

MACRO aor221d4
    CLASS CORE ;
    FOREIGN aor221d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.530 2.920 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.270 2.020 2.180 2.460 ;
        RECT  1.270 2.020 1.510 2.920 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.700 2.740 3.580 ;
        RECT  1.870 2.700 2.740 2.940 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.500 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.890 3.140 4.420 3.580 ;
        RECT  3.890 2.500 4.150 3.580 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.987  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.850 3.190 6.570 3.590 ;
        RECT  6.330 1.640 6.570 3.590 ;
        RECT  6.170 1.640 6.570 2.050 ;
        RECT  4.870 1.640 6.570 1.880 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.600 4.620 6.000 5.600 ;
        RECT  4.330 4.190 4.570 5.600 ;
        RECT  2.850 4.300 3.090 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.660 0.000 5.900 1.270 ;
        RECT  4.140 0.000 4.380 1.270 ;
        RECT  2.230 0.000 2.470 1.300 ;
        RECT  0.260 0.000 0.500 1.780 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.730 4.080 1.130 4.620 ;
        RECT  0.730 4.380 2.470 4.620 ;
        RECT  1.470 3.610 1.870 4.060 ;
        RECT  1.470 3.820 3.910 4.060 ;
        RECT  0.770 1.540 4.630 1.780 ;
        RECT  4.390 1.540 4.630 2.900 ;
        RECT  4.390 2.500 5.500 2.900 ;
        RECT  0.770 1.540 1.010 3.410 ;
        RECT  0.150 3.170 1.010 3.410 ;
    END
END aor221d4

MACRO aor221d2
    CLASS CORE ;
    FOREIGN aor221d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.530 2.920 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.270 2.020 2.180 2.460 ;
        RECT  1.270 2.020 1.510 3.040 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.720 2.740 3.580 ;
        RECT  1.950 2.720 2.740 2.960 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.500 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.850 3.140 4.420 3.580 ;
        RECT  3.850 2.500 4.090 3.580 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.370  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.870 3.190 5.540 3.590 ;
        RECT  5.300 1.540 5.540 3.590 ;
        RECT  4.910 1.540 5.540 1.790 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.690 4.180 5.930 5.600 ;
        RECT  4.340 4.190 4.580 5.600 ;
        RECT  2.840 4.300 3.080 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.690 0.000 5.930 1.270 ;
        RECT  4.340 0.000 4.580 1.270 ;
        RECT  2.230 0.000 2.470 1.300 ;
        RECT  0.260 0.000 0.500 1.780 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.730 4.200 1.130 4.620 ;
        RECT  0.730 4.380 2.440 4.620 ;
        RECT  1.470 3.610 1.870 4.060 ;
        RECT  1.470 3.820 3.920 4.060 ;
        RECT  0.770 1.540 4.590 1.780 ;
        RECT  4.350 1.540 4.590 2.900 ;
        RECT  4.350 2.500 4.850 2.900 ;
        RECT  0.770 1.540 1.010 3.490 ;
        RECT  0.150 3.250 1.010 3.490 ;
    END
END aor221d2

MACRO aor221d1
    CLASS CORE ;
    FOREIGN aor221d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.530 2.920 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.270 2.020 2.180 2.460 ;
        RECT  1.270 2.020 1.510 3.040 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.720 2.740 3.580 ;
        RECT  1.950 2.720 2.740 2.960 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.020 3.500 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 3.140 4.420 3.580 ;
        RECT  3.980 2.500 4.220 3.580 ;
        RECT  3.770 2.500 4.220 2.900 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.214  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.860 3.100 5.480 3.500 ;
        RECT  5.100 1.460 5.480 3.500 ;
        RECT  5.050 1.460 5.480 1.860 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.340 4.190 4.580 5.600 ;
        RECT  2.840 4.300 3.080 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.340 0.000 4.580 1.270 ;
        RECT  2.230 0.000 2.470 1.300 ;
        RECT  0.260 0.000 0.500 1.780 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.730 4.200 1.130 4.620 ;
        RECT  0.730 4.380 2.440 4.620 ;
        RECT  1.470 3.610 1.870 4.060 ;
        RECT  1.470 3.820 3.920 4.060 ;
        RECT  0.770 1.540 4.770 1.780 ;
        RECT  4.510 1.540 4.770 2.390 ;
        RECT  0.770 1.540 1.010 3.490 ;
        RECT  0.150 3.250 1.010 3.490 ;
    END
END aor221d1

MACRO aor21d4
    CLASS CORE ;
    FOREIGN aor21d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.500 2.560 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.580 2.220 2.180 2.460 ;
        RECT  1.740 2.020 2.180 2.460 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.580 3.300 3.020 ;
        RECT  2.420 2.580 3.300 2.900 ;
        RECT  2.420 2.500 2.820 2.900 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.131  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.750 3.130 5.450 3.450 ;
        RECT  4.940 3.040 5.450 3.450 ;
        RECT  4.940 1.460 5.340 3.450 ;
        RECT  4.540 1.460 5.340 1.900 ;
        RECT  3.610 1.460 5.340 1.700 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.280 4.620 4.680 5.600 ;
        RECT  2.980 4.620 3.380 5.600 ;
        RECT  1.710 4.710 2.110 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.350 0.000 4.750 0.980 ;
        RECT  2.840 0.000 3.240 0.890 ;
        RECT  0.410 0.000 0.650 1.140 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.890 3.260 2.840 3.500 ;
        RECT  1.120 3.310 2.200 3.550 ;
        RECT  1.340 1.380 1.740 1.780 ;
        RECT  0.740 1.540 3.370 1.780 ;
        RECT  3.130 1.540 3.370 2.340 ;
        RECT  3.130 2.100 3.760 2.340 ;
        RECT  0.740 1.540 0.980 3.110 ;
        RECT  0.410 2.870 0.780 3.550 ;
    END
END aor21d4

MACRO aor21d2
    CLASS CORE ;
    FOREIGN aor21d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.460 2.500 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.490 1.640 3.020 ;
        RECT  1.400 2.100 1.640 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.420  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.090 2.020 2.740 2.500 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.256  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.360 3.140 3.860 3.940 ;
        RECT  3.530 1.020 3.770 3.940 ;
        RECT  3.160 1.020 3.770 1.300 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  4.010 4.430 4.250 5.600 ;
        RECT  2.590 4.710 2.990 5.600 ;
        RECT  1.500 4.710 1.900 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  4.010 0.000 4.250 1.420 ;
        RECT  2.440 0.000 2.680 1.300 ;
        RECT  0.270 0.000 0.510 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.170 3.050 2.410 4.030 ;
        RECT  0.730 3.790 2.410 4.030 ;
        RECT  0.700 1.540 3.220 1.780 ;
        RECT  0.700 1.540 1.150 1.970 ;
        RECT  2.980 1.540 3.220 2.500 ;
        RECT  0.700 1.540 0.940 3.370 ;
        RECT  0.150 3.130 0.940 3.370 ;
    END
END aor21d2

MACRO aor21d1
    CLASS CORE ;
    FOREIGN aor21d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.460 2.500 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.490 1.640 3.020 ;
        RECT  1.400 2.100 1.640 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.420  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.090 2.020 2.740 2.500 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.034  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.370 3.140 3.800 3.940 ;
        RECT  3.560 1.020 3.800 3.940 ;
        RECT  3.370 1.020 3.800 1.340 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  2.760 4.710 3.170 5.600 ;
        RECT  1.500 4.710 1.900 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  2.440 0.000 2.680 1.300 ;
        RECT  0.270 0.000 0.510 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.180 3.050 2.420 4.030 ;
        RECT  0.730 3.790 2.420 4.030 ;
        RECT  0.700 1.540 3.220 1.780 ;
        RECT  0.700 1.540 1.150 1.970 ;
        RECT  2.980 1.540 3.220 2.500 ;
        RECT  0.700 1.540 0.940 3.370 ;
        RECT  0.150 3.130 0.940 3.370 ;
    END
END aor21d1

MACRO aor211d4
    CLASS CORE ;
    FOREIGN aor211d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.497  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.470 0.500 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.477  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 3.700 1.620 4.140 ;
        RECT  1.220 2.470 1.620 2.870 ;
        RECT  1.220 2.470 1.460 4.140 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.415  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.970 2.320 2.740 2.560 ;
        RECT  2.300 2.020 2.740 2.560 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.429  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  2.980 2.580 3.860 2.900 ;
        RECT  2.980 2.500 3.380 2.900 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.131  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.310 3.130 6.010 3.450 ;
        RECT  5.500 3.040 6.010 3.450 ;
        RECT  5.500 1.460 5.900 3.450 ;
        RECT  5.100 1.460 5.900 1.900 ;
        RECT  4.170 1.460 5.900 1.700 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.840 4.620 5.240 5.600 ;
        RECT  3.540 4.620 3.940 5.600 ;
        RECT  2.370 3.890 2.610 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.910 0.000 5.310 0.980 ;
        RECT  3.400 0.000 3.800 0.890 ;
        RECT  0.900 0.000 1.140 1.370 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.700 3.130 2.600 3.370 ;
        RECT  2.360 3.260 3.400 3.500 ;
        RECT  1.580 1.540 3.930 1.780 ;
        RECT  0.150 1.660 2.040 1.900 ;
        RECT  0.150 1.660 0.980 1.930 ;
        RECT  1.800 1.540 2.040 1.980 ;
        RECT  3.690 1.540 3.930 2.340 ;
        RECT  3.690 2.100 4.320 2.340 ;
        RECT  0.740 1.660 0.980 3.560 ;
        RECT  0.270 3.320 0.980 3.560 ;
    END
END aor211d4

MACRO aor211d2
    CLASS CORE ;
    FOREIGN aor211d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.515  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.020 0.500 2.870 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.499  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.700 1.460 3.940 ;
        RECT  1.220 2.470 1.460 3.940 ;
        RECT  0.620 3.700 1.060 4.140 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.250 2.540 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.449  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  3.420 3.010 3.660 4.140 ;
        RECT  2.260 3.010 3.660 3.250 ;
        RECT  2.260 2.850 2.660 3.250 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.234  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.580 4.420 3.450 ;
        RECT  4.180 1.670 4.420 3.450 ;
        RECT  3.750 1.670 4.420 1.910 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.570 4.120 4.810 5.600 ;
        RECT  3.120 4.410 3.520 5.600 ;
        RECT  2.210 4.410 2.610 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.490 0.000 4.890 1.420 ;
        RECT  2.780 0.000 3.180 1.300 ;
        RECT  0.790 0.000 1.190 1.140 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.700 3.580 2.970 3.820 ;
        RECT  1.700 3.580 1.940 4.500 ;
        RECT  1.270 4.260 1.940 4.500 ;
        RECT  1.560 1.380 1.960 1.780 ;
        RECT  0.150 1.540 3.200 1.780 ;
        RECT  2.960 1.540 3.200 2.440 ;
        RECT  2.960 2.200 3.660 2.440 ;
        RECT  0.740 1.540 0.980 3.370 ;
        RECT  0.150 3.130 0.980 3.370 ;
    END
END aor211d2

MACRO aor211d1
    CLASS CORE ;
    FOREIGN aor211d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.460 2.920 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.496  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 1.620 2.550 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.220 3.580 ;
        RECT  1.980 2.520 2.220 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.570 3.300 3.580 ;
        RECT  2.580 2.570 3.300 2.810 ;
        END
    END C2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.005  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.930 3.150 4.360 3.550 ;
        RECT  4.110 1.560 4.360 3.550 ;
        RECT  4.010 1.560 4.360 2.530 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.440 3.890 3.680 5.600 ;
        RECT  1.810 4.710 2.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.020 0.000 3.260 1.300 ;
        RECT  0.830 0.000 1.070 1.140 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.230 4.020 3.060 4.260 ;
        RECT  0.150 1.540 3.770 1.780 ;
        RECT  3.530 1.540 3.770 2.500 ;
        RECT  0.700 1.540 0.940 3.400 ;
        RECT  0.150 3.160 0.940 3.400 ;
    END
END aor211d1

MACRO aon211d4
    CLASS CORE ;
    FOREIGN aon211d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.660 2.750 3.020 ;
        RECT  2.430 2.450 2.750 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.020 2.180 2.380 ;
        RECT  1.770 2.020 2.010 2.710 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.460 0.460 2.500 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.478  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.310 3.580 ;
        RECT  1.070 2.290 1.310 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.113  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.800 3.500 6.570 3.740 ;
        RECT  4.860 1.840 6.570 2.080 ;
        RECT  5.660 1.840 6.100 3.740 ;
        RECT  4.860 1.840 6.100 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.540 4.620 5.940 5.600 ;
        RECT  4.190 4.710 4.590 5.600 ;
        RECT  2.820 4.710 3.220 5.600 ;
        RECT  0.970 4.440 1.210 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.680 0.000 5.920 1.280 ;
        RECT  4.350 0.000 4.590 1.280 ;
        RECT  2.100 0.000 2.500 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.570 3.060 1.810 4.060 ;
        RECT  0.150 3.820 1.810 4.060 ;
        RECT  0.150 0.980 1.260 1.220 ;
        RECT  1.020 0.980 1.260 1.510 ;
        RECT  1.020 1.270 2.460 1.510 ;
        RECT  2.780 1.760 3.240 2.170 ;
        RECT  3.000 2.380 4.100 2.620 ;
        RECT  3.000 1.760 3.240 3.500 ;
        RECT  2.230 3.260 3.240 3.500 ;
        RECT  3.500 1.850 4.590 2.090 ;
        RECT  4.350 2.440 5.160 2.680 ;
        RECT  4.350 1.850 4.590 3.370 ;
        RECT  3.500 3.130 4.590 3.370 ;
    END
END aon211d4

MACRO aon211d2
    CLASS CORE ;
    FOREIGN aon211d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 2.440 2.750 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.020 2.100 2.460 ;
        RECT  1.770 2.020 2.010 2.920 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.460 0.460 2.500 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.479  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.310 3.580 ;
        RECT  1.070 2.290 1.310 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.513  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.930 3.130 5.520 3.450 ;
        RECT  5.280 1.770 5.520 3.450 ;
        RECT  5.100 2.580 5.520 3.450 ;
        RECT  4.870 1.770 5.520 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.550 4.710 5.950 5.600 ;
        RECT  4.190 4.710 4.590 5.600 ;
        RECT  2.840 4.710 3.240 5.600 ;
        RECT  0.990 4.300 1.230 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.690 0.000 5.930 1.360 ;
        RECT  4.360 0.000 4.600 1.360 ;
        RECT  2.150 0.000 2.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.580 3.360 1.820 4.060 ;
        RECT  0.150 3.820 1.820 4.060 ;
        RECT  0.150 0.980 1.760 1.220 ;
        RECT  1.520 0.980 1.760 1.510 ;
        RECT  1.520 1.270 2.460 1.510 ;
        RECT  2.800 1.770 3.240 2.170 ;
        RECT  3.000 2.380 4.110 2.620 ;
        RECT  3.000 1.770 3.240 3.500 ;
        RECT  2.240 3.260 3.240 3.500 ;
        RECT  3.510 1.850 4.590 2.090 ;
        RECT  4.350 2.360 4.860 2.760 ;
        RECT  4.350 1.850 4.590 3.370 ;
        RECT  3.510 3.130 4.590 3.370 ;
    END
END aon211d2

MACRO aon211d1
    CLASS CORE ;
    FOREIGN aon211d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.494  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 2.580 2.750 3.020 ;
        RECT  2.510 2.350 2.750 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.940 2.180 2.440 ;
        RECT  1.770 1.940 2.010 2.820 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.487  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.020 0.460 2.960 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.310 3.580 ;
        RECT  1.070 2.320 1.310 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.202  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.240 3.260 3.240 3.500 ;
        RECT  3.000 1.460 3.240 3.500 ;
        RECT  2.860 1.460 3.240 2.130 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.890 4.130 3.130 5.600 ;
        RECT  0.990 4.300 1.230 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  1.070 0.000 1.470 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.580 3.060 1.820 4.060 ;
        RECT  0.150 3.820 1.820 4.060 ;
        RECT  2.140 1.160 2.460 1.500 ;
        RECT  0.150 1.260 2.460 1.500 ;
    END
END aon211d1

MACRO aoim3m11d4
    CLASS CORE ;
    FOREIGN aoim3m11d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.554  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.920 3.700 5.540 4.140 ;
        RECT  4.920 2.190 5.480 2.430 ;
        RECT  4.920 2.190 5.160 4.140 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.413  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.070 3.580 ;
        RECT  0.620 2.540 0.860 3.580 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.493  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 1.720 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.516  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.360 3.580 ;
        RECT  2.120 2.230 2.360 3.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.441  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.080 3.160 3.860 3.580 ;
        RECT  3.080 2.670 3.360 3.580 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.997  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.210 3.290 9.920 3.530 ;
        RECT  8.210 1.850 9.920 2.090 ;
        RECT  9.020 1.850 9.460 3.530 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  8.860 4.340 9.100 5.600 ;
        RECT  7.550 4.340 7.790 5.600 ;
        RECT  3.640 4.590 4.040 5.600 ;
        RECT  0.300 4.700 0.700 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  9.030 0.000 9.270 1.310 ;
        RECT  7.720 0.000 7.960 1.310 ;
        RECT  5.690 0.000 5.930 1.340 ;
        RECT  4.390 0.000 4.630 1.340 ;
        RECT  2.170 0.000 2.570 0.980 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.570 1.300 3.310 1.540 ;
        RECT  3.070 1.300 3.310 2.430 ;
        RECT  2.600 2.190 4.040 2.430 ;
        RECT  2.600 2.190 2.840 4.140 ;
        RECT  1.610 3.900 2.840 4.140 ;
        RECT  0.120 1.240 0.550 1.640 ;
        RECT  0.120 1.240 0.360 4.190 ;
        RECT  0.120 3.870 1.330 4.190 ;
        RECT  4.360 2.670 4.600 4.210 ;
        RECT  3.080 3.970 4.600 4.210 ;
        RECT  1.090 3.870 1.330 4.620 ;
        RECT  3.080 3.970 3.320 4.620 ;
        RECT  1.090 4.380 3.320 4.620 ;
        RECT  3.570 1.020 4.150 1.270 ;
        RECT  3.910 1.020 4.150 1.900 ;
        RECT  3.910 1.660 6.040 1.900 ;
        RECT  5.800 2.600 7.490 2.840 ;
        RECT  5.800 1.660 6.040 3.460 ;
        RECT  5.480 3.200 6.040 3.460 ;
        RECT  6.870 1.850 7.970 2.090 ;
        RECT  7.730 2.600 8.520 2.840 ;
        RECT  7.730 1.850 7.970 3.530 ;
        RECT  6.870 3.290 7.970 3.530 ;
    END
END aoim3m11d4

MACRO aoim3m11d2
    CLASS CORE ;
    FOREIGN aoim3m11d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.560  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.920 2.580 5.540 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.413  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.070 3.580 ;
        RECT  0.620 2.540 0.860 3.580 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.493  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.890 1.620 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.516  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.190 3.580 ;
        RECT  1.950 2.390 2.190 3.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.441  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.080 3.140 3.860 3.580 ;
        RECT  3.080 2.670 3.320 3.580 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.370  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.260 3.130 7.410 3.370 ;
        RECT  6.260 1.460 7.320 1.980 ;
        RECT  6.260 1.460 6.500 3.370 ;
        RECT  6.220 1.460 7.320 1.900 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.890 4.180 8.130 5.600 ;
        RECT  6.520 4.180 6.760 5.600 ;
        RECT  3.450 4.710 3.850 5.600 ;
        RECT  0.300 4.710 0.700 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.660 0.000 7.900 1.340 ;
        RECT  5.690 0.000 5.930 1.340 ;
        RECT  4.390 0.000 4.630 1.340 ;
        RECT  2.170 0.000 2.570 0.980 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.570 1.300 3.310 1.540 ;
        RECT  3.070 1.300 3.310 2.430 ;
        RECT  2.450 2.190 4.040 2.430 ;
        RECT  2.450 2.190 2.690 4.140 ;
        RECT  1.610 3.900 2.690 4.140 ;
        RECT  0.120 1.240 0.550 1.640 ;
        RECT  4.100 2.670 4.680 3.070 ;
        RECT  0.120 1.240 0.360 4.190 ;
        RECT  0.120 3.870 1.370 4.190 ;
        RECT  1.130 3.870 1.370 4.620 ;
        RECT  2.950 4.220 4.340 4.460 ;
        RECT  4.100 2.670 4.340 4.460 ;
        RECT  1.130 4.380 3.190 4.620 ;
        RECT  3.570 1.020 4.150 1.270 ;
        RECT  3.910 1.020 4.150 1.900 ;
        RECT  3.910 1.660 5.950 1.900 ;
        RECT  5.710 1.660 5.950 2.330 ;
        RECT  8.120 2.290 8.360 3.250 ;
        RECT  7.680 3.010 8.360 3.250 ;
        RECT  5.210 3.280 6.020 3.520 ;
        RECT  5.780 2.090 6.020 3.930 ;
        RECT  7.680 3.010 7.920 3.930 ;
        RECT  5.780 3.690 7.920 3.930 ;
        RECT  7.570 1.580 8.840 1.900 ;
        RECT  7.570 1.580 7.810 2.460 ;
        RECT  7.030 2.220 7.810 2.460 ;
        RECT  8.600 1.580 8.840 3.920 ;
        RECT  8.410 3.510 8.840 3.920 ;
    END
END aoim3m11d2

MACRO aoim3m11d1
    CLASS CORE ;
    FOREIGN aoim3m11d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.536  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.920 3.700 5.540 4.140 ;
        RECT  4.920 2.190 5.480 2.430 ;
        RECT  4.920 2.190 5.160 4.140 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.413  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.070 3.580 ;
        RECT  0.620 2.540 0.860 3.580 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.493  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 1.720 2.460 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.516  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.360 3.580 ;
        RECT  2.120 2.230 2.360 3.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.441  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.080 3.160 3.860 3.580 ;
        RECT  3.080 2.670 3.360 3.580 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.650  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.420 3.200 6.040 3.460 ;
        RECT  5.800 1.660 6.040 3.460 ;
        RECT  5.720 1.660 6.040 2.460 ;
        RECT  3.910 1.660 6.040 1.900 ;
        RECT  3.910 1.020 4.150 1.900 ;
        RECT  3.570 1.020 4.150 1.270 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  3.560 4.590 3.960 5.600 ;
        RECT  0.450 4.710 0.850 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.690 0.000 5.930 1.340 ;
        RECT  4.390 0.000 4.630 1.340 ;
        RECT  2.170 0.000 2.570 0.980 ;
        RECT  0.740 0.000 1.140 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.570 1.300 3.310 1.540 ;
        RECT  3.070 1.300 3.310 2.430 ;
        RECT  2.600 2.190 4.040 2.430 ;
        RECT  2.600 2.190 2.840 4.140 ;
        RECT  1.560 3.900 2.840 4.140 ;
        RECT  0.120 1.240 0.550 1.640 ;
        RECT  0.120 1.240 0.360 4.310 ;
        RECT  0.120 3.790 0.470 4.310 ;
        RECT  4.360 2.670 4.600 4.210 ;
        RECT  3.080 3.970 4.600 4.210 ;
        RECT  0.120 4.070 1.320 4.310 ;
        RECT  1.080 4.070 1.320 4.620 ;
        RECT  3.080 3.970 3.320 4.620 ;
        RECT  1.080 4.380 3.320 4.620 ;
    END
END aoim3m11d1

MACRO aoim31d4
    CLASS CORE ;
    FOREIGN aoim31d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.040 2.340 3.290 3.100 ;
        RECT  2.940 3.100 3.280 3.580 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.503  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.460 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.300 1.610 3.020 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 3.140 2.180 3.580 ;
        RECT  1.860 2.390 2.100 3.580 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.997  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.410 3.290 7.120 3.530 ;
        RECT  5.410 1.850 7.120 2.090 ;
        RECT  6.220 1.850 6.660 3.530 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.060 4.340 6.300 5.600 ;
        RECT  4.750 4.340 4.990 5.600 ;
        RECT  1.990 4.480 2.230 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.230 0.000 6.470 1.310 ;
        RECT  4.920 0.000 5.160 1.310 ;
        RECT  3.450 0.000 3.690 1.470 ;
        RECT  2.120 0.000 2.360 1.470 ;
        RECT  0.800 0.000 1.040 1.470 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.700 1.820 1.860 2.060 ;
        RECT  0.150 1.850 0.940 2.090 ;
        RECT  0.700 1.820 0.940 4.160 ;
        RECT  2.460 3.040 2.700 4.160 ;
        RECT  0.150 3.920 2.700 4.160 ;
        RECT  2.780 1.850 3.800 2.090 ;
        RECT  3.560 2.600 4.690 2.840 ;
        RECT  3.560 1.850 3.800 4.500 ;
        RECT  3.370 4.100 3.800 4.500 ;
        RECT  4.070 1.850 5.170 2.090 ;
        RECT  4.930 2.600 5.720 2.840 ;
        RECT  4.930 1.850 5.170 3.380 ;
        RECT  4.070 3.140 5.170 3.380 ;
    END
END aoim31d4

MACRO aoim31d2
    CLASS CORE ;
    FOREIGN aoim31d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.040 2.340 3.290 3.100 ;
        RECT  2.940 3.100 3.280 3.580 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.503  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.460 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.300 1.610 3.020 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 3.140 2.180 3.580 ;
        RECT  1.860 2.390 2.100 3.580 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.263  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.410 3.290 6.200 3.530 ;
        RECT  5.960 1.770 6.200 3.530 ;
        RECT  5.660 1.770 6.200 2.460 ;
        RECT  5.410 1.770 6.200 2.170 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  6.060 4.340 6.300 5.600 ;
        RECT  4.750 4.340 4.990 5.600 ;
        RECT  1.990 4.480 2.230 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  6.230 0.000 6.470 1.480 ;
        RECT  4.920 0.000 5.160 1.480 ;
        RECT  3.450 0.000 3.690 1.470 ;
        RECT  2.120 0.000 2.360 1.470 ;
        RECT  0.800 0.000 1.040 1.470 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.700 1.820 1.860 2.060 ;
        RECT  0.150 1.850 0.940 2.090 ;
        RECT  0.700 1.820 0.940 4.160 ;
        RECT  2.460 3.040 2.700 4.160 ;
        RECT  0.150 3.920 2.700 4.160 ;
        RECT  2.780 1.850 3.800 2.090 ;
        RECT  3.560 2.600 4.690 2.840 ;
        RECT  3.560 1.850 3.800 4.500 ;
        RECT  3.370 4.100 3.800 4.500 ;
        RECT  4.070 1.850 5.170 2.090 ;
        RECT  4.930 2.720 5.720 2.960 ;
        RECT  4.930 1.850 5.170 3.530 ;
        RECT  4.070 3.290 5.170 3.530 ;
    END
END aoim31d2

MACRO aoim31d1
    CLASS CORE ;
    FOREIGN aoim31d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.040 2.340 3.290 3.100 ;
        RECT  2.940 3.100 3.280 3.580 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.503  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.460 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.300 1.610 3.020 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 3.140 2.180 3.580 ;
        RECT  1.860 2.390 2.100 3.580 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.363  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.370 4.100 3.800 4.500 ;
        RECT  3.560 1.850 3.800 4.500 ;
        RECT  3.490 3.700 3.800 4.500 ;
        RECT  2.780 1.850 3.800 2.090 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  1.990 4.480 2.230 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  3.450 0.000 3.690 1.470 ;
        RECT  2.120 0.000 2.360 1.470 ;
        RECT  0.800 0.000 1.040 1.470 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.700 1.820 1.860 2.060 ;
        RECT  0.150 1.850 0.940 2.090 ;
        RECT  0.700 1.820 0.940 4.160 ;
        RECT  2.460 3.040 2.700 4.160 ;
        RECT  0.150 3.920 2.700 4.160 ;
    END
END aoim31d1

MACRO aoim311d4
    CLASS CORE ;
    FOREIGN aoim311d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.575  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.110 2.580 4.980 3.010 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.540  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 3.700 3.340 4.140 ;
        RECT  3.100 2.640 3.340 4.140 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.447  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.460 2.950 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.230 3.580 ;
        RECT  0.980 2.670 1.230 3.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.650 2.540 2.180 3.020 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.097  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.350 1.460 6.660 1.810 ;
        RECT  4.820 3.260 6.530 3.500 ;
        RECT  5.350 1.460 6.250 1.900 ;
        RECT  5.350 1.460 5.590 3.500 ;
        RECT  4.940 1.460 6.660 1.800 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  6.750 4.620 7.150 5.600 ;
        RECT  5.360 4.620 5.760 5.600 ;
        RECT  2.090 4.610 2.490 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  6.990 0.000 7.400 0.980 ;
        RECT  5.670 0.000 6.080 0.980 ;
        RECT  3.750 0.000 3.990 1.420 ;
        RECT  2.330 0.000 2.570 1.420 ;
        RECT  0.970 0.000 1.210 1.280 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 1.870 1.780 ;
        RECT  1.470 1.700 2.660 1.940 ;
        RECT  2.420 1.700 2.660 3.500 ;
        RECT  2.210 3.260 2.450 4.110 ;
        RECT  0.150 3.870 2.450 4.110 ;
        RECT  2.930 1.850 4.640 2.090 ;
        RECT  3.630 1.850 3.870 4.360 ;
        RECT  7.270 2.520 7.510 4.360 ;
        RECT  3.630 4.120 7.510 4.360 ;
        RECT  7.740 1.480 7.990 2.280 ;
        RECT  6.750 2.040 7.990 2.280 ;
        RECT  6.750 2.040 6.990 2.890 ;
        RECT  5.880 2.490 6.990 2.890 ;
        RECT  7.750 1.480 7.990 3.450 ;
    END
END aoim311d4

MACRO aoim311d2
    CLASS CORE ;
    FOREIGN aoim311d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.400 2.020 4.980 2.460 ;
        RECT  4.400 2.020 4.640 2.860 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.520 3.590 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.000 0.490 2.920 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 2.520 1.620 2.920 ;
        RECT  0.620 3.720 1.450 4.140 ;
        RECT  1.210 2.520 1.450 4.140 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.220 3.580 ;
        RECT  1.980 2.520 2.220 3.580 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.333  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.140 5.790 3.580 ;
        RECT  5.230 1.410 5.780 1.730 ;
        RECT  5.230 1.410 5.470 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.220 4.300 6.460 5.600 ;
        RECT  4.900 4.300 5.140 5.600 ;
        RECT  2.230 3.870 2.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.120 0.000 6.520 0.980 ;
        RECT  4.820 0.000 5.220 0.980 ;
        RECT  3.480 0.000 3.880 0.980 ;
        RECT  1.550 0.000 1.790 1.590 ;
        RECT  0.230 0.000 0.470 1.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.730 1.750 1.130 2.150 ;
        RECT  0.730 1.830 3.140 2.150 ;
        RECT  0.730 1.750 0.970 3.410 ;
        RECT  0.270 3.170 0.970 3.410 ;
        RECT  2.820 0.990 3.060 1.560 ;
        RECT  2.820 1.320 4.070 1.560 ;
        RECT  3.830 1.470 4.480 1.710 ;
        RECT  3.830 1.320 4.070 3.370 ;
        RECT  6.400 2.520 6.640 3.300 ;
        RECT  3.830 3.130 4.860 3.370 ;
        RECT  4.620 3.130 4.860 4.060 ;
        RECT  6.240 3.060 6.480 4.060 ;
        RECT  4.620 3.820 6.480 4.060 ;
        RECT  6.780 1.410 7.020 2.260 ;
        RECT  5.710 2.020 7.160 2.260 ;
        RECT  6.920 2.020 7.160 3.940 ;
        RECT  6.720 3.540 7.160 3.940 ;
    END
END aoim311d2

MACRO aoim311d1
    CLASS CORE ;
    FOREIGN aoim311d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.530 2.020 5.000 2.820 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.553  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 3.140 3.710 3.580 ;
        RECT  3.470 2.220 3.710 3.580 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.940 0.630 2.340 ;
        RECT  0.120 1.450 0.480 2.340 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.370 3.020 ;
        RECT  0.970 1.980 1.370 3.020 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.610 2.020 2.180 2.460 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.928  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.020 1.340 4.740 1.580 ;
        RECT  3.950 3.130 4.720 3.450 ;
        RECT  3.950 1.340 4.190 3.450 ;
        RECT  3.420 1.340 4.190 1.880 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  2.220 4.600 2.620 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.920 0.000 5.320 0.980 ;
        RECT  3.600 0.000 4.000 0.980 ;
        RECT  1.460 0.000 1.860 0.980 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 1.340 2.660 1.580 ;
        RECT  2.230 1.340 2.660 1.740 ;
        RECT  2.420 2.070 3.110 2.310 ;
        RECT  2.420 1.340 2.660 2.940 ;
        RECT  2.380 2.700 2.620 3.500 ;
        RECT  0.250 3.260 2.620 3.500 ;
    END
END aoim311d1

MACRO aoim2m11d4
    CLASS CORE ;
    FOREIGN aoim2m11d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 3.120 4.440 3.580 ;
        RECT  4.200 2.750 4.440 3.580 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.442  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.540 1.060 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 2.310 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.260 3.020 ;
        RECT  1.860 2.210 2.260 3.020 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.018  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.530 3.290 8.240 3.530 ;
        RECT  6.530 1.850 8.240 2.090 ;
        RECT  7.340 1.850 7.780 3.530 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.180 4.340 7.420 5.600 ;
        RECT  5.870 4.340 6.110 5.600 ;
        RECT  2.610 4.460 2.850 5.600 ;
        RECT  0.800 4.360 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.350 0.000 7.590 1.280 ;
        RECT  6.040 0.000 6.280 1.280 ;
        RECT  3.930 0.000 4.170 1.420 ;
        RECT  2.520 0.000 2.760 1.220 ;
        RECT  0.970 0.000 1.210 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.630 0.980 2.280 1.220 ;
        RECT  2.040 0.980 2.280 1.700 ;
        RECT  2.040 1.460 2.790 1.700 ;
        RECT  2.550 2.730 3.230 2.970 ;
        RECT  2.550 1.460 2.790 3.600 ;
        RECT  1.420 3.360 2.790 3.600 ;
        RECT  0.120 1.380 0.550 1.780 ;
        RECT  3.500 2.150 3.920 2.470 ;
        RECT  0.120 1.380 0.360 4.120 ;
        RECT  0.120 3.530 0.550 4.120 ;
        RECT  3.500 2.150 3.740 4.120 ;
        RECT  0.120 3.870 3.740 4.120 ;
        RECT  3.110 1.670 4.920 1.910 ;
        RECT  4.480 1.620 4.920 2.020 ;
        RECT  4.680 2.600 5.810 2.840 ;
        RECT  4.680 1.620 4.920 4.220 ;
        RECT  4.490 3.820 4.920 4.220 ;
        RECT  5.190 1.850 6.290 2.090 ;
        RECT  6.050 2.600 6.840 2.840 ;
        RECT  6.050 1.850 6.290 3.530 ;
        RECT  5.190 3.290 6.290 3.530 ;
    END
END aoim2m11d4

MACRO aoim2m11d2
    CLASS CORE ;
    FOREIGN aoim2m11d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 3.120 4.440 3.580 ;
        RECT  4.200 2.750 4.440 3.580 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.442  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.540 1.060 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 2.310 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.260 3.020 ;
        RECT  1.860 2.210 2.260 3.020 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.263  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.530 3.290 7.320 3.530 ;
        RECT  7.080 1.770 7.320 3.530 ;
        RECT  6.780 1.770 7.320 2.460 ;
        RECT  6.530 1.770 7.320 2.170 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  7.180 4.340 7.420 5.600 ;
        RECT  5.870 4.340 6.110 5.600 ;
        RECT  2.610 4.460 2.850 5.600 ;
        RECT  0.800 4.360 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  7.350 0.000 7.590 1.480 ;
        RECT  6.040 0.000 6.280 1.480 ;
        RECT  3.930 0.000 4.170 1.420 ;
        RECT  2.520 0.000 2.760 1.220 ;
        RECT  0.970 0.000 1.210 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.630 0.980 2.280 1.220 ;
        RECT  2.040 0.980 2.280 1.700 ;
        RECT  2.040 1.460 2.790 1.700 ;
        RECT  2.550 2.730 3.230 2.970 ;
        RECT  2.550 1.460 2.790 3.600 ;
        RECT  1.420 3.360 2.790 3.600 ;
        RECT  0.120 1.380 0.550 1.780 ;
        RECT  3.500 2.150 3.920 2.470 ;
        RECT  0.120 1.380 0.360 4.120 ;
        RECT  0.120 3.530 0.550 4.120 ;
        RECT  3.500 2.150 3.740 4.120 ;
        RECT  0.120 3.870 3.740 4.120 ;
        RECT  3.110 1.670 4.920 1.910 ;
        RECT  4.480 1.620 4.920 2.020 ;
        RECT  4.680 2.600 5.810 2.840 ;
        RECT  4.680 1.620 4.920 4.220 ;
        RECT  4.490 3.820 4.920 4.220 ;
        RECT  5.190 1.850 6.290 2.090 ;
        RECT  6.050 2.720 6.840 2.960 ;
        RECT  6.050 1.850 6.290 3.530 ;
        RECT  5.190 3.290 6.290 3.530 ;
    END
END aoim2m11d2

MACRO aoim2m11d1
    CLASS CORE ;
    FOREIGN aoim2m11d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 3.120 4.440 3.580 ;
        RECT  4.200 2.750 4.440 3.580 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.442  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.540 1.060 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 2.310 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.260 3.020 ;
        RECT  1.860 2.210 2.260 3.020 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.749  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.490 3.820 4.920 4.220 ;
        RECT  4.680 1.620 4.920 4.220 ;
        RECT  4.600 1.620 4.920 2.460 ;
        RECT  4.480 1.620 4.920 2.020 ;
        RECT  3.110 1.670 4.920 1.910 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  2.610 4.460 2.850 5.600 ;
        RECT  0.800 4.360 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.930 0.000 4.170 1.420 ;
        RECT  2.520 0.000 2.760 1.220 ;
        RECT  0.970 0.000 1.210 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.630 0.980 2.280 1.220 ;
        RECT  2.040 0.980 2.280 1.700 ;
        RECT  2.040 1.460 2.790 1.700 ;
        RECT  2.550 2.730 3.230 2.970 ;
        RECT  2.550 1.460 2.790 3.600 ;
        RECT  1.420 3.360 2.790 3.600 ;
        RECT  0.120 1.380 0.550 1.780 ;
        RECT  3.500 2.150 3.920 2.470 ;
        RECT  0.120 1.380 0.360 4.120 ;
        RECT  0.120 3.530 0.550 4.120 ;
        RECT  3.500 2.150 3.740 4.120 ;
        RECT  0.120 3.870 3.740 4.120 ;
    END
END aoim2m11d1

MACRO aoim22d4
    CLASS CORE ;
    FOREIGN aoim22d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.369  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.540 2.890 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.369  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.480 3.580 ;
        RECT  1.100 2.970 1.480 3.580 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.506  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.190 2.580 3.860 3.040 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.506  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.540 2.740 3.450 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.215  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.380 1.600 6.020 1.840 ;
        RECT  4.280 3.900 6.010 4.140 ;
        RECT  5.100 3.700 5.550 4.140 ;
        RECT  5.310 1.600 5.550 4.140 ;
        RECT  4.380 1.600 5.550 1.850 ;
        RECT  4.380 1.270 4.620 1.850 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.030 4.620 5.430 5.600 ;
        RECT  3.420 4.610 3.820 5.600 ;
        RECT  1.660 4.610 2.060 5.600 ;
        RECT  0.230 4.080 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.120 0.000 5.360 1.100 ;
        RECT  3.610 0.000 4.010 0.980 ;
        RECT  1.180 0.000 1.580 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.310 1.960 1.550 ;
        RECT  1.720 1.700 3.660 1.940 ;
        RECT  3.420 1.700 3.660 2.320 ;
        RECT  1.540 2.290 1.960 2.690 ;
        RECT  1.720 1.310 1.960 4.060 ;
        RECT  0.890 3.820 1.960 4.060 ;
        RECT  2.400 1.220 4.140 1.460 ;
        RECT  3.900 1.220 4.140 2.330 ;
        RECT  4.120 2.090 4.360 3.660 ;
        RECT  3.570 3.420 4.360 3.660 ;
        RECT  3.570 3.420 3.810 4.090 ;
        RECT  2.260 3.850 3.810 4.090 ;
    END
END aoim22d4

MACRO aoim22d2
    CLASS CORE ;
    FOREIGN aoim22d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.540 2.890 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.380 3.580 ;
        RECT  1.140 2.690 1.380 3.580 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.487  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.340 2.570 3.860 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.487  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.580 2.860 3.440 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.266  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.290 3.740 4.980 4.140 ;
        RECT  4.540 3.700 4.980 4.140 ;
        RECT  4.640 1.390 4.880 4.140 ;
        RECT  4.480 1.390 4.880 1.790 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.940 4.510 5.180 5.600 ;
        RECT  3.500 4.510 3.740 5.600 ;
        RECT  1.660 4.510 2.060 5.600 ;
        RECT  0.230 4.080 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  5.110 0.000 5.350 1.100 ;
        RECT  3.610 0.000 4.010 0.980 ;
        RECT  1.180 0.000 1.580 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.310 2.060 1.550 ;
        RECT  1.820 2.000 3.760 2.240 ;
        RECT  1.820 1.310 2.060 4.060 ;
        RECT  0.890 3.820 2.060 4.060 ;
        RECT  2.400 1.420 4.240 1.660 ;
        RECT  4.000 1.420 4.240 2.350 ;
        RECT  4.120 2.110 4.360 3.500 ;
        RECT  3.650 3.260 4.360 3.500 ;
        RECT  3.650 3.260 3.890 3.930 ;
        RECT  2.320 3.690 3.890 3.930 ;
    END
END aoim22d2

MACRO aoim22d1
    CLASS CORE ;
    FOREIGN aoim22d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.650  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.460 3.300 1.900 ;
        RECT  2.600 2.580 3.220 2.820 ;
        RECT  2.980 1.460 3.220 2.820 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.649  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.460 2.180 3.800 3.580 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.347  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.540 2.890 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.347  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.820 2.300 1.400 2.540 ;
        RECT  1.160 1.820 1.400 2.540 ;
        RECT  0.620 3.140 1.060 3.580 ;
        RECT  0.820 2.300 1.060 3.580 ;
        END
    END B2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.543  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.120 3.140 3.060 3.580 ;
        RECT  2.350 1.650 2.590 2.340 ;
        RECT  2.120 2.100 2.360 3.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  1.380 4.510 1.780 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  3.340 0.000 3.770 0.980 ;
        RECT  1.470 0.000 1.870 0.890 ;
        RECT  0.230 0.000 0.470 1.630 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 1.310 1.880 1.550 ;
        RECT  1.640 1.310 1.880 3.690 ;
        RECT  1.380 3.450 1.880 3.690 ;
        RECT  1.380 3.450 1.620 4.080 ;
        RECT  0.150 3.840 1.620 4.080 ;
        RECT  1.990 3.910 3.770 4.150 ;
    END
END aoim22d1

MACRO aoim21d4
    CLASS CORE ;
    FOREIGN aoim21d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.459  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.440 2.520 2.680 3.580 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.460 2.400 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.240 3.020 ;
        RECT  1.000 2.130 1.240 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.997  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.850 3.290 6.560 3.530 ;
        RECT  4.850 1.850 6.560 2.090 ;
        RECT  5.660 1.850 6.100 3.530 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.500 4.340 5.740 5.600 ;
        RECT  4.190 4.340 4.430 5.600 ;
        RECT  1.440 3.890 1.680 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.670 0.000 5.910 1.310 ;
        RECT  4.360 0.000 4.600 1.310 ;
        RECT  2.890 0.000 3.130 1.480 ;
        RECT  1.540 0.000 1.780 1.410 ;
        RECT  0.230 0.000 0.470 1.210 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 1.470 1.120 1.890 ;
        RECT  0.720 1.650 1.820 1.890 ;
        RECT  1.580 2.520 2.060 2.920 ;
        RECT  1.580 1.650 1.820 3.500 ;
        RECT  0.150 3.260 1.820 3.500 ;
        RECT  2.060 1.730 3.240 1.970 ;
        RECT  3.000 2.600 4.130 2.840 ;
        RECT  3.000 1.730 3.240 4.060 ;
        RECT  2.610 3.820 3.240 4.060 ;
        RECT  3.510 1.850 4.610 2.090 ;
        RECT  4.370 2.600 5.160 2.840 ;
        RECT  4.370 1.850 4.610 3.530 ;
        RECT  3.510 3.290 4.610 3.530 ;
    END
END aoim21d4

MACRO aoim21d2
    CLASS CORE ;
    FOREIGN aoim21d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.459  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.440 2.520 2.680 3.580 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.460 2.400 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.240 3.020 ;
        RECT  1.000 2.130 1.240 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.263  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.850 3.290 5.640 3.530 ;
        RECT  5.400 1.770 5.640 3.530 ;
        RECT  5.100 1.770 5.640 2.460 ;
        RECT  4.850 1.770 5.640 2.170 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.500 4.340 5.740 5.600 ;
        RECT  4.190 4.340 4.430 5.600 ;
        RECT  1.440 3.890 1.680 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.670 0.000 5.910 1.480 ;
        RECT  4.360 0.000 4.600 1.480 ;
        RECT  2.890 0.000 3.130 1.480 ;
        RECT  1.540 0.000 1.780 1.410 ;
        RECT  0.230 0.000 0.470 1.210 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 1.470 1.120 1.890 ;
        RECT  0.720 1.650 1.820 1.890 ;
        RECT  1.580 2.520 2.060 2.920 ;
        RECT  1.580 1.650 1.820 3.500 ;
        RECT  0.150 3.260 1.820 3.500 ;
        RECT  2.060 1.730 3.240 1.970 ;
        RECT  3.000 2.600 4.130 2.840 ;
        RECT  3.000 1.730 3.240 4.060 ;
        RECT  2.610 3.820 3.240 4.060 ;
        RECT  3.510 1.850 4.610 2.090 ;
        RECT  4.370 2.720 5.160 2.960 ;
        RECT  4.370 1.850 4.610 3.530 ;
        RECT  3.510 3.290 4.610 3.530 ;
    END
END aoim21d2

MACRO aoim21d1
    CLASS CORE ;
    FOREIGN aoim21d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.459  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.740 3.580 ;
        RECT  2.440 2.520 2.680 3.580 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.460 2.400 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.240 3.020 ;
        RECT  1.000 2.130 1.240 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.385  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.610 3.820 3.240 4.060 ;
        RECT  3.000 1.730 3.240 4.060 ;
        RECT  2.920 1.730 3.240 2.460 ;
        RECT  2.060 1.730 3.240 1.970 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  1.440 3.890 1.680 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.890 0.000 3.130 1.480 ;
        RECT  1.540 0.000 1.780 1.410 ;
        RECT  0.230 0.000 0.470 1.210 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 1.470 1.120 1.890 ;
        RECT  0.720 1.650 1.820 1.890 ;
        RECT  1.580 2.520 2.060 2.920 ;
        RECT  1.580 1.650 1.820 3.500 ;
        RECT  0.150 3.260 1.820 3.500 ;
    END
END aoim21d1

MACRO aoim211d4
    CLASS CORE ;
    FOREIGN aoim211d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.499  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.300 3.300 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.700 2.740 4.140 ;
        RECT  2.380 2.590 2.620 4.140 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.471  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.460 2.960 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.230 3.580 ;
        RECT  0.990 2.660 1.230 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.997  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.410 3.290 7.120 3.530 ;
        RECT  5.410 1.850 7.120 2.090 ;
        RECT  6.220 1.850 6.660 3.530 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.060 4.340 6.300 5.600 ;
        RECT  4.750 4.340 4.990 5.600 ;
        RECT  1.520 4.300 1.760 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.230 0.000 6.470 1.310 ;
        RECT  4.920 0.000 5.160 1.310 ;
        RECT  2.880 0.000 3.120 1.400 ;
        RECT  1.540 0.000 1.780 1.310 ;
        RECT  0.230 0.000 0.470 1.310 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 1.670 1.780 1.910 ;
        RECT  1.540 2.600 2.000 2.990 ;
        RECT  1.540 1.670 1.780 4.060 ;
        RECT  0.150 3.820 1.780 4.060 ;
        RECT  0.150 3.820 0.550 4.400 ;
        RECT  2.050 1.670 3.780 1.930 ;
        RECT  3.370 1.670 3.780 2.070 ;
        RECT  3.540 2.600 4.690 2.840 ;
        RECT  3.540 1.670 3.780 3.800 ;
        RECT  3.270 3.380 3.780 3.800 ;
        RECT  4.070 1.850 5.170 2.090 ;
        RECT  4.930 2.600 5.720 2.840 ;
        RECT  4.930 1.850 5.170 3.530 ;
        RECT  4.070 3.290 5.170 3.530 ;
    END
END aoim211d4

MACRO aoim211d2
    CLASS CORE ;
    FOREIGN aoim211d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.499  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.300 3.300 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.467  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.700 2.740 4.140 ;
        RECT  2.380 2.590 2.620 4.140 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.471  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.460 2.960 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.230 3.580 ;
        RECT  0.990 2.660 1.230 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.263  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.410 3.290 6.200 3.530 ;
        RECT  5.960 1.770 6.200 3.530 ;
        RECT  5.660 1.770 6.200 2.460 ;
        RECT  5.410 1.770 6.200 2.170 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  6.060 4.340 6.300 5.600 ;
        RECT  4.750 4.340 4.990 5.600 ;
        RECT  1.520 4.300 1.760 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  6.230 0.000 6.470 1.480 ;
        RECT  4.920 0.000 5.160 1.480 ;
        RECT  2.880 0.000 3.120 1.400 ;
        RECT  1.540 0.000 1.780 1.310 ;
        RECT  0.230 0.000 0.470 1.310 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 1.670 1.780 1.910 ;
        RECT  1.540 2.600 2.000 2.990 ;
        RECT  1.540 1.670 1.780 4.060 ;
        RECT  0.150 3.820 1.780 4.060 ;
        RECT  0.150 3.820 0.550 4.400 ;
        RECT  2.050 1.670 3.780 1.930 ;
        RECT  3.370 1.670 3.780 2.070 ;
        RECT  3.540 2.600 4.690 2.840 ;
        RECT  3.540 1.670 3.780 3.800 ;
        RECT  3.270 3.380 3.780 3.800 ;
        RECT  4.070 1.850 5.170 2.090 ;
        RECT  4.930 2.720 5.720 2.960 ;
        RECT  4.930 1.850 5.170 3.530 ;
        RECT  4.070 3.290 5.170 3.530 ;
    END
END aoim211d2

MACRO aoim211d1
    CLASS CORE ;
    FOREIGN aoim211d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.499  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.320 3.300 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.700 2.740 4.140 ;
        RECT  2.380 2.590 2.620 4.140 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.471  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.460 2.960 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.230 3.580 ;
        RECT  0.990 2.660 1.230 3.580 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.603  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.270 3.300 3.780 4.140 ;
        RECT  3.540 1.690 3.780 4.140 ;
        RECT  3.370 1.690 3.780 2.090 ;
        RECT  2.050 1.690 3.780 1.950 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  1.520 4.300 1.760 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  2.880 0.000 3.120 1.420 ;
        RECT  1.540 0.000 1.780 1.330 ;
        RECT  0.230 0.000 0.470 1.330 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 1.690 1.780 1.930 ;
        RECT  1.540 2.600 2.000 2.990 ;
        RECT  1.540 1.690 1.780 4.060 ;
        RECT  0.150 3.820 1.780 4.060 ;
        RECT  0.150 3.820 0.550 4.400 ;
    END
END aoim211d1

MACRO aoi322d4
    CLASS CORE ;
    FOREIGN aoi322d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.421  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.520 1.320 3.050 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.442  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.540 2.170 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 1.970 2.740 2.670 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.110 2.020 3.860 2.460 ;
        RECT  2.970 2.840 3.370 3.240 ;
        RECT  3.110 2.020 3.370 3.240 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.410 3.700 6.100 4.140 ;
        RECT  5.410 2.680 5.650 4.140 ;
        RECT  5.220 2.680 5.650 3.080 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.509  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.460 2.180 4.980 2.580 ;
        RECT  4.550 2.020 4.980 2.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.990 2.860 4.420 3.580 ;
        RECT  3.720 2.700 4.120 3.100 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.122  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.250 3.050 8.810 3.580 ;
        RECT  8.410 1.220 8.810 3.580 ;
        RECT  7.100 1.220 8.810 1.460 ;
        RECT  7.100 1.000 7.500 1.460 ;
        RECT  7.090 4.020 7.490 4.420 ;
        RECT  7.250 3.050 7.490 4.420 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.830 4.550 8.230 5.600 ;
        RECT  6.350 4.550 6.750 5.600 ;
        RECT  5.390 4.440 5.790 5.600 ;
        RECT  4.090 4.440 4.490 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.840 0.000 8.240 0.980 ;
        RECT  6.440 0.000 6.680 1.420 ;
        RECT  3.220 0.000 3.620 0.980 ;
        RECT  0.460 0.000 0.700 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 4.260 3.190 4.500 ;
        RECT  2.040 3.480 3.750 3.880 ;
        RECT  3.350 3.820 5.050 4.060 ;
        RECT  1.560 1.180 2.010 1.620 ;
        RECT  1.560 1.220 5.340 1.620 ;
        RECT  4.880 1.580 5.650 1.750 ;
        RECT  5.150 1.580 5.650 1.850 ;
        RECT  5.410 1.580 5.650 2.380 ;
        RECT  5.410 2.140 6.400 2.380 ;
        RECT  5.990 2.140 6.400 2.760 ;
        RECT  1.560 1.180 1.800 3.610 ;
        RECT  0.720 3.360 1.800 3.610 ;
        RECT  5.580 1.100 6.130 1.340 ;
        RECT  5.890 1.100 6.130 1.900 ;
        RECT  5.890 1.660 6.880 1.900 ;
        RECT  6.640 2.360 7.960 2.760 ;
        RECT  6.640 1.660 6.880 3.370 ;
        RECT  5.920 3.130 6.880 3.370 ;
    END
END aoi322d4

MACRO aoi322d2
    CLASS CORE ;
    FOREIGN aoi322d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.421  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.550 1.330 3.050 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.442  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.540 2.170 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 1.970 2.740 2.800 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.120 2.020 3.860 2.460 ;
        RECT  2.980 2.710 3.380 3.110 ;
        RECT  3.120 2.020 3.380 3.110 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.410 3.700 6.100 4.140 ;
        RECT  5.410 2.680 5.650 4.140 ;
        RECT  5.220 2.680 5.650 3.080 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.509  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.460 2.180 4.980 2.580 ;
        RECT  4.550 2.020 4.980 2.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 2.840 4.420 3.580 ;
        RECT  3.720 2.700 4.120 3.100 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.230 3.050 7.860 3.580 ;
        RECT  7.620 1.220 7.860 3.580 ;
        RECT  7.110 1.220 7.860 1.460 ;
        RECT  7.110 1.000 7.510 1.460 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.870 4.140 8.110 5.600 ;
        RECT  6.570 3.720 6.810 5.600 ;
        RECT  5.470 4.440 5.710 5.600 ;
        RECT  4.170 4.440 4.410 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.850 0.000 8.250 0.980 ;
        RECT  6.400 0.000 6.640 1.420 ;
        RECT  3.220 0.000 3.620 0.980 ;
        RECT  0.460 0.000 0.700 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 4.380 3.190 4.620 ;
        RECT  2.050 3.670 3.750 3.940 ;
        RECT  3.350 3.820 5.050 4.060 ;
        RECT  1.570 1.180 2.010 1.620 ;
        RECT  1.570 1.220 5.340 1.620 ;
        RECT  4.880 1.580 5.650 1.750 ;
        RECT  5.150 1.580 5.650 1.850 ;
        RECT  5.410 1.580 5.650 2.380 ;
        RECT  5.410 2.140 6.400 2.380 ;
        RECT  5.990 2.140 6.400 2.580 ;
        RECT  1.570 1.180 1.810 3.950 ;
        RECT  0.710 3.700 1.810 3.950 ;
        RECT  5.580 1.100 6.130 1.340 ;
        RECT  5.890 1.100 6.130 1.900 ;
        RECT  5.890 1.660 6.880 1.900 ;
        RECT  6.640 2.020 7.380 2.420 ;
        RECT  6.640 1.660 6.880 3.370 ;
        RECT  5.920 3.130 6.880 3.370 ;
    END
END aoi322d2

MACRO aoi322d1
    CLASS CORE ;
    FOREIGN aoi322d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.421  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.520 1.320 3.050 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.442  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.460 0.540 2.170 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 2.580 2.740 3.240 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.970 3.860 2.460 ;
        RECT  2.860 1.970 3.860 2.370 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 3.080 5.650 3.580 ;
        RECT  5.220 2.680 5.650 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.509  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.400 2.180 4.980 2.580 ;
        RECT  4.550 2.020 4.980 2.580 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.488  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.990 2.860 4.420 3.580 ;
        RECT  3.720 2.700 4.120 3.100 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.729  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.730 1.220 5.130 1.620 ;
        RECT  1.560 1.220 5.130 1.540 ;
        RECT  1.560 1.220 2.180 1.900 ;
        RECT  0.720 3.360 1.800 3.610 ;
        RECT  1.560 1.220 1.800 3.610 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.390 4.440 5.790 5.600 ;
        RECT  4.090 4.440 4.490 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  3.070 0.000 3.470 0.980 ;
        RECT  0.460 0.000 0.700 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 4.260 3.190 4.500 ;
        RECT  2.040 3.480 3.750 3.880 ;
        RECT  3.350 3.820 5.050 4.060 ;
    END
END aoi322d1

MACRO aoi321d4
    CLASS CORE ;
    FOREIGN aoi321d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.352  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.490 0.550 2.900 ;
        RECT  0.120 2.010 0.500 2.900 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.130 2.740 3.580 ;
        RECT  1.670 2.820 2.540 3.220 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.350 2.460 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.479  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.520 2.870 4.980 3.610 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.840 2.380 4.240 2.900 ;
        RECT  2.860 2.380 4.240 2.620 ;
        RECT  2.860 2.020 3.300 2.620 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.479  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.100 3.140 3.860 3.580 ;
        RECT  3.100 2.860 3.500 3.580 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.133  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.540 4.050 8.250 4.290 ;
        RECT  8.010 1.460 8.250 4.290 ;
        RECT  7.850 3.050 8.250 4.290 ;
        RECT  6.550 1.460 8.250 1.900 ;
        RECT  6.540 4.050 6.940 4.450 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.270 4.530 7.680 5.600 ;
        RECT  5.800 4.470 6.210 5.600 ;
        RECT  4.590 4.540 4.990 5.600 ;
        RECT  3.290 4.540 3.690 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.130 0.000 7.530 1.150 ;
        RECT  5.790 0.000 6.190 1.170 ;
        RECT  2.200 0.000 2.600 0.890 ;
        RECT  0.230 0.000 0.470 1.620 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 4.180 1.120 4.620 ;
        RECT  0.720 4.380 2.390 4.620 ;
        RECT  1.420 3.580 1.820 4.110 ;
        RECT  1.420 3.870 4.430 4.110 ;
        RECT  0.820 1.380 4.960 1.780 ;
        RECT  4.720 1.380 4.960 2.630 ;
        RECT  4.720 2.390 5.830 2.630 ;
        RECT  5.430 2.390 5.830 2.810 ;
        RECT  0.820 1.380 1.060 3.670 ;
        RECT  0.150 3.430 1.060 3.670 ;
        RECT  5.220 1.570 6.310 1.810 ;
        RECT  6.070 2.420 7.230 2.800 ;
        RECT  6.070 1.570 6.310 3.370 ;
        RECT  5.330 3.130 6.310 3.370 ;
    END
END aoi321d4

MACRO aoi321d2
    CLASS CORE ;
    FOREIGN aoi321d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.352  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.490 0.550 2.900 ;
        RECT  0.120 2.010 0.500 2.900 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.130 2.740 3.580 ;
        RECT  1.670 2.820 2.540 3.220 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.350 2.460 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.479  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.520 2.870 4.980 3.610 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.840 2.380 4.240 2.900 ;
        RECT  2.860 2.380 4.240 2.620 ;
        RECT  2.860 2.020 3.300 2.620 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.479  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.100 3.140 3.860 3.580 ;
        RECT  3.100 2.860 3.500 3.580 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.483  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.660 3.130 7.280 3.370 ;
        RECT  7.040 1.460 7.280 3.370 ;
        RECT  6.660 1.460 7.280 1.900 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  7.240 4.410 7.650 5.600 ;
        RECT  5.910 4.460 6.320 5.600 ;
        RECT  4.590 4.540 4.990 5.600 ;
        RECT  3.290 4.540 3.690 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  7.240 0.000 7.640 1.150 ;
        RECT  5.900 0.000 6.300 1.170 ;
        RECT  2.200 0.000 2.600 0.890 ;
        RECT  0.230 0.000 0.470 1.620 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 4.180 1.120 4.620 ;
        RECT  0.720 4.380 2.390 4.620 ;
        RECT  1.420 3.580 1.820 4.110 ;
        RECT  1.420 3.870 4.430 4.110 ;
        RECT  0.820 1.380 5.040 1.780 ;
        RECT  4.800 1.380 5.040 2.630 ;
        RECT  4.800 2.390 5.940 2.630 ;
        RECT  5.540 2.390 5.940 2.810 ;
        RECT  0.820 1.380 1.060 3.670 ;
        RECT  0.150 3.430 1.060 3.670 ;
        RECT  5.330 1.570 6.420 1.810 ;
        RECT  6.180 2.420 6.800 2.800 ;
        RECT  6.180 1.570 6.420 3.370 ;
        RECT  5.330 3.130 6.420 3.370 ;
    END
END aoi321d2

MACRO aoi321d1
    CLASS CORE ;
    FOREIGN aoi321d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.352  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.490 0.550 2.900 ;
        RECT  0.120 2.010 0.500 2.900 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.130 2.740 3.580 ;
        RECT  1.670 2.820 2.540 3.220 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.020 2.350 2.460 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.479  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 1.920 4.980 2.490 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.840 2.380 4.240 2.900 ;
        RECT  2.860 2.380 4.240 2.620 ;
        RECT  2.860 2.020 3.300 2.620 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.479  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.100 3.140 3.860 3.580 ;
        RECT  3.100 2.860 3.500 3.580 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.491  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.130 4.800 1.370 ;
        RECT  0.820 1.130 1.230 1.610 ;
        RECT  0.150 3.430 1.060 3.670 ;
        RECT  0.820 1.130 1.060 3.670 ;
        RECT  0.620 3.130 1.060 3.670 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.590 4.540 4.990 5.600 ;
        RECT  3.290 4.540 3.690 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  2.200 0.000 2.600 0.890 ;
        RECT  0.230 0.000 0.470 1.620 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 4.180 1.120 4.620 ;
        RECT  0.720 4.380 2.390 4.620 ;
        RECT  1.420 3.580 1.820 4.110 ;
        RECT  1.420 3.870 4.430 4.110 ;
    END
END aoi321d1

MACRO aoi31d4
    CLASS CORE ;
    FOREIGN aoi31d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.350 2.250 2.810 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.250 2.110 3.580 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.460 1.620 1.910 ;
        RECT  1.080 2.250 1.480 2.650 ;
        RECT  1.180 1.460 1.480 2.650 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.500 0.800 2.900 ;
        RECT  0.120 2.020 0.500 2.900 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.975  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.860 1.770 6.570 2.170 ;
        RECT  4.830 3.140 6.540 3.610 ;
        RECT  5.840 1.770 6.080 3.610 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.570 4.170 5.970 5.600 ;
        RECT  4.270 4.620 4.670 5.600 ;
        RECT  1.310 4.710 1.710 5.600 ;
        RECT  0.150 3.160 0.550 3.560 ;
        RECT  0.150 3.160 0.390 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.600 0.000 6.000 1.260 ;
        RECT  4.300 0.000 4.700 1.260 ;
        RECT  2.630 0.000 3.030 1.430 ;
        RECT  0.150 0.000 0.550 1.430 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 3.970 2.480 4.210 ;
        RECT  2.030 1.770 3.290 2.010 ;
        RECT  3.050 2.450 3.520 2.850 ;
        RECT  3.050 1.770 3.290 3.660 ;
        RECT  2.710 3.260 3.290 3.660 ;
        RECT  3.530 1.750 4.000 2.170 ;
        RECT  3.760 2.450 5.520 2.850 ;
        RECT  3.760 1.750 4.000 3.490 ;
        RECT  3.530 3.090 4.000 3.490 ;
    END
END aoi31d4

MACRO aoi31d2
    CLASS CORE ;
    FOREIGN aoi31d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.431  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.220 0.460 3.030 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.530 1.620 3.100 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.860 2.250 2.280 2.650 ;
        RECT  1.860 1.460 2.180 2.650 ;
        RECT  1.740 1.460 2.180 1.910 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.550 2.550 3.300 3.040 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.313  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 4.020 4.140 ;
        RECT  3.560 3.460 4.020 4.140 ;
        RECT  3.560 1.720 4.020 2.120 ;
        RECT  3.560 1.720 3.800 4.140 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.180 4.340 4.580 5.600 ;
        RECT  2.800 4.630 3.200 5.600 ;
        RECT  2.880 3.340 3.120 5.600 ;
        RECT  1.560 3.340 3.120 3.580 ;
        RECT  0.330 4.790 0.730 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.280 0.000 4.680 0.940 ;
        RECT  2.920 0.000 3.320 0.940 ;
        RECT  0.150 0.000 0.550 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.890 3.970 2.640 4.210 ;
        RECT  0.890 0.980 2.680 1.220 ;
        RECT  2.440 0.980 2.680 1.480 ;
        RECT  2.440 1.240 4.810 1.480 ;
        RECT  4.570 1.240 4.810 2.420 ;
        RECT  0.890 0.980 1.130 2.100 ;
        RECT  4.570 2.020 5.000 2.420 ;
        RECT  0.700 1.680 0.940 3.640 ;
        RECT  0.150 3.340 0.940 3.640 ;
        RECT  0.150 3.340 0.550 3.740 ;
        RECT  5.050 1.330 5.480 1.750 ;
        RECT  4.040 2.690 4.440 3.110 ;
        RECT  4.040 2.850 5.480 3.110 ;
        RECT  5.240 1.330 5.480 3.640 ;
        RECT  4.970 2.850 5.480 3.640 ;
    END
END aoi31d2

MACRO aoi31d1
    CLASS CORE ;
    FOREIGN aoi31d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.420  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.220 0.460 3.030 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.414  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.530 1.630 3.100 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.414  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.720 2.280 2.650 ;
        RECT  1.740 1.460 2.180 1.910 ;
        END
    END B2
    PIN B3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.700 2.620 3.240 3.040 ;
        RECT  2.860 1.930 3.240 3.040 ;
        END
    END B3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.065  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.460 1.130 2.100 ;
        RECT  0.150 3.340 0.940 3.640 ;
        RECT  0.700 1.460 0.940 3.640 ;
        RECT  0.620 1.460 1.130 1.900 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.800 4.630 3.200 5.600 ;
        RECT  2.880 3.340 3.120 5.600 ;
        RECT  1.560 3.340 3.120 3.580 ;
        RECT  0.330 4.790 0.730 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.830 0.000 3.180 1.520 ;
        RECT  0.150 0.000 0.550 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.890 3.970 2.640 4.210 ;
    END
END aoi31d1

MACRO aoi311d4
    CLASS CORE ;
    FOREIGN aoi311d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 3.140 1.060 3.580 ;
        RECT  0.600 2.170 0.920 3.580 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.750 1.700 2.150 ;
        RECT  1.180 1.750 1.620 2.460 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.130 2.180 3.580 ;
        RECT  1.840 2.960 2.180 3.580 ;
        RECT  1.840 2.560 2.160 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.499  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.430 2.020 3.300 2.460 ;
        RECT  2.430 2.020 2.850 2.770 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.530 2.550 3.930 2.950 ;
        RECT  3.420 3.140 3.860 3.580 ;
        RECT  3.530 2.550 3.860 3.580 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.217  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.730 3.130 7.160 4.600 ;
        RECT  6.780 1.460 7.160 4.600 ;
        RECT  6.720 1.460 7.160 1.930 ;
        RECT  5.420 3.130 7.160 3.370 ;
        RECT  5.420 1.460 7.160 1.900 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  5.980 4.410 6.380 5.600 ;
        RECT  4.640 4.580 5.050 5.600 ;
        RECT  3.490 4.700 3.890 5.600 ;
        RECT  2.100 4.300 2.500 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  5.980 0.000 6.400 1.150 ;
        RECT  4.660 0.000 5.080 1.170 ;
        RECT  3.400 0.000 3.800 0.980 ;
        RECT  1.110 0.000 1.510 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.740 3.270 3.090 4.060 ;
        RECT  1.350 3.820 3.090 4.060 ;
        RECT  1.350 3.820 1.770 4.430 ;
        RECT  0.120 1.090 0.550 1.510 ;
        RECT  0.120 1.270 3.780 1.510 ;
        RECT  3.540 1.270 3.780 2.300 ;
        RECT  3.540 2.060 4.700 2.300 ;
        RECT  4.290 2.060 4.700 2.340 ;
        RECT  0.120 1.090 0.360 4.250 ;
        RECT  0.120 3.850 0.560 4.250 ;
        RECT  4.100 1.570 5.180 1.810 ;
        RECT  4.940 2.200 6.110 2.440 ;
        RECT  4.940 1.570 5.180 3.370 ;
        RECT  4.100 3.130 5.180 3.370 ;
    END
END aoi311d4

MACRO aoi311d2
    CLASS CORE ;
    FOREIGN aoi311d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 3.140 1.060 3.580 ;
        RECT  0.600 2.170 0.920 3.580 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.750 1.700 2.150 ;
        RECT  1.180 1.750 1.620 2.460 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.840 2.560 2.190 2.960 ;
        RECT  1.740 3.130 2.180 3.580 ;
        RECT  1.840 2.560 2.180 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.510 2.020 3.300 2.460 ;
        RECT  2.510 2.020 2.910 2.770 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.560 2.550 3.970 2.960 ;
        RECT  3.420 3.140 3.860 3.580 ;
        RECT  3.560 2.550 3.860 3.580 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.530  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.500 3.130 6.100 3.370 ;
        RECT  5.860 1.460 6.100 3.370 ;
        RECT  5.500 1.460 6.100 1.900 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  6.060 4.410 6.470 5.600 ;
        RECT  4.720 4.410 5.140 5.600 ;
        RECT  3.490 4.700 3.900 5.600 ;
        RECT  2.160 4.300 2.560 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  6.070 0.000 6.470 1.150 ;
        RECT  4.730 0.000 5.130 1.170 ;
        RECT  3.460 0.000 3.860 0.980 ;
        RECT  1.110 0.000 1.510 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.720 3.310 3.120 4.060 ;
        RECT  1.400 3.820 3.120 4.060 ;
        RECT  1.400 3.820 1.820 4.430 ;
        RECT  0.120 1.090 0.550 1.510 ;
        RECT  0.120 1.270 3.920 1.510 ;
        RECT  3.680 1.270 3.920 2.300 ;
        RECT  3.680 2.060 4.780 2.300 ;
        RECT  4.380 2.060 4.780 2.340 ;
        RECT  0.120 1.090 0.360 4.250 ;
        RECT  0.120 3.850 0.560 4.250 ;
        RECT  4.160 1.570 5.260 1.810 ;
        RECT  5.020 2.200 5.620 2.440 ;
        RECT  5.020 1.570 5.260 3.370 ;
        RECT  4.150 3.130 5.260 3.370 ;
    END
END aoi311d2

MACRO aoi311d1
    CLASS CORE ;
    FOREIGN aoi311d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.210 1.010 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.523  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.300 2.200 1.720 2.600 ;
        RECT  1.220 3.140 1.620 3.580 ;
        RECT  1.300 2.200 1.620 3.580 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.527  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.000 2.160 2.680 2.560 ;
        RECT  2.350 1.450 2.680 2.560 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.548  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.920 2.020 3.300 2.460 ;
        RECT  2.530 2.840 3.160 3.240 ;
        RECT  2.920 2.020 3.160 3.240 ;
        END
    END C2
    PIN C3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.568  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.840 3.800 4.140 ;
        END
    END C3
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.654  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.660 2.110 1.900 ;
        RECT  1.710 1.410 2.110 1.900 ;
        RECT  0.140 1.490 0.560 1.900 ;
        RECT  0.140 3.250 0.550 3.650 ;
        RECT  0.140 3.250 0.500 4.140 ;
        RECT  0.140 1.490 0.380 4.140 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  3.370 4.620 3.770 5.600 ;
        RECT  2.040 4.620 2.440 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  3.370 0.000 3.770 0.980 ;
        RECT  0.890 0.000 1.290 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.780 3.810 3.180 4.380 ;
        RECT  1.300 4.140 3.180 4.380 ;
        RECT  1.300 4.140 1.700 4.540 ;
    END
END aoi311d1

MACRO aoi22d4
    CLASS CORE ;
    FOREIGN aoi22d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.460 2.130 2.640 ;
        RECT  0.620 1.460 2.130 1.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.870 2.020 3.300 2.810 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.110 2.570 1.620 3.020 ;
        RECT  1.110 2.240 1.510 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.494  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.170 0.790 2.570 ;
        RECT  0.120 2.170 0.500 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.161  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.860 3.050 6.570 3.450 ;
        RECT  4.860 1.460 6.570 1.900 ;
        RECT  5.300 1.460 5.580 3.450 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.600 4.040 6.000 5.600 ;
        RECT  4.300 4.430 4.700 5.600 ;
        RECT  0.800 4.080 1.200 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.600 0.000 6.000 0.980 ;
        RECT  4.300 0.000 4.700 0.980 ;
        RECT  2.890 0.000 3.130 1.490 ;
        RECT  0.150 0.000 0.550 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.390 1.850 3.630 ;
        RECT  1.450 3.390 1.850 4.400 ;
        RECT  1.440 4.160 3.210 4.400 ;
        RECT  1.530 0.980 2.630 1.220 ;
        RECT  3.840 2.520 4.080 3.450 ;
        RECT  2.180 3.210 4.080 3.450 ;
        RECT  2.390 0.980 2.630 3.580 ;
        RECT  2.180 3.140 2.630 3.580 ;
        RECT  3.510 1.540 4.560 1.780 ;
        RECT  4.320 2.390 5.020 2.790 ;
        RECT  4.320 1.540 4.560 3.930 ;
        RECT  3.510 3.690 4.560 3.930 ;
    END
END aoi22d4

MACRO aoi22d2
    CLASS CORE ;
    FOREIGN aoi22d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.460 2.130 2.640 ;
        RECT  0.620 1.460 2.130 1.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.870 2.020 3.300 2.810 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.110 2.570 1.620 3.020 ;
        RECT  1.110 2.240 1.510 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.494  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.170 0.790 2.570 ;
        RECT  0.120 2.170 0.500 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.517  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.990 3.050 5.580 3.450 ;
        RECT  5.300 1.380 5.580 3.450 ;
        RECT  4.870 1.380 5.580 1.900 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.600 4.000 6.000 5.600 ;
        RECT  4.250 4.430 4.650 5.600 ;
        RECT  0.800 4.080 1.200 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.610 0.000 6.010 0.980 ;
        RECT  4.310 0.000 4.710 0.980 ;
        RECT  2.890 0.000 3.130 1.490 ;
        RECT  0.150 0.000 0.550 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.390 1.850 3.630 ;
        RECT  1.450 3.390 1.850 4.400 ;
        RECT  1.440 4.160 3.210 4.400 ;
        RECT  1.530 0.980 2.630 1.220 ;
        RECT  3.840 2.520 4.080 3.450 ;
        RECT  2.180 3.210 4.080 3.450 ;
        RECT  2.390 0.980 2.630 3.580 ;
        RECT  2.180 3.140 2.630 3.580 ;
        RECT  3.510 1.540 4.560 1.780 ;
        RECT  4.320 2.140 5.020 2.540 ;
        RECT  4.320 1.540 4.560 3.930 ;
        RECT  3.510 3.690 4.560 3.930 ;
    END
END aoi22d2

MACRO aoi22d1
    CLASS CORE ;
    FOREIGN aoi22d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.230 1.460 2.740 1.900 ;
        RECT  1.230 1.460 1.470 2.640 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.490 2.810 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.570 2.250 3.020 ;
        RECT  1.850 2.240 2.250 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.494  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.170 3.240 3.020 ;
        RECT  2.570 2.170 3.240 2.570 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.572  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.980 1.830 1.220 ;
        RECT  0.620 3.140 1.180 3.580 ;
        RECT  0.730 0.980 0.970 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.160 4.430 2.560 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.890 0.000 3.130 1.220 ;
        RECT  0.230 0.000 0.470 1.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.510 3.390 3.210 3.630 ;
        RECT  1.510 3.390 1.910 4.400 ;
        RECT  0.150 4.160 1.920 4.400 ;
    END
END aoi22d1

MACRO aoi222d4
    CLASS CORE ;
    FOREIGN aoi222d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.310 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.910 0.800 2.310 ;
        RECT  0.120 1.460 0.500 2.310 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.670 2.000 2.070 ;
        RECT  1.180 1.460 1.620 2.070 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.700 2.720 2.460 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.506  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.440 2.520 4.040 2.920 ;
        RECT  3.440 2.020 3.860 2.920 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.527  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.340 2.020 4.980 2.700 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.419  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.390 1.770 7.510 2.170 ;
        RECT  5.390 3.310 7.100 3.710 ;
        RECT  5.390 3.140 6.100 3.710 ;
        RECT  5.390 1.770 5.630 3.710 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.270 4.450 7.670 5.600 ;
        RECT  5.960 4.450 6.360 5.600 ;
        RECT  4.070 4.340 4.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.820 0.000 8.220 0.980 ;
        RECT  6.370 0.000 6.770 0.980 ;
        RECT  4.780 0.000 5.180 0.980 ;
        RECT  2.690 0.000 3.090 0.980 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 4.260 3.170 4.500 ;
        RECT  2.030 3.560 5.030 3.800 ;
        RECT  1.350 0.980 2.450 1.220 ;
        RECT  2.210 1.220 7.990 1.460 ;
        RECT  7.750 1.220 7.990 2.460 ;
        RECT  7.750 2.060 8.150 2.460 ;
        RECT  2.960 1.220 3.200 2.940 ;
        RECT  1.550 2.700 3.200 2.940 ;
        RECT  1.550 2.700 1.790 3.500 ;
        RECT  0.720 3.260 1.790 3.500 ;
        RECT  0.720 3.260 1.120 4.020 ;
        RECT  0.720 3.780 1.130 4.020 ;
        RECT  8.390 1.430 8.790 1.820 ;
        RECT  6.410 2.440 7.350 2.940 ;
        RECT  6.410 2.700 8.630 2.940 ;
        RECT  8.390 1.430 8.630 3.450 ;
        RECT  8.000 2.700 8.630 3.450 ;
    END
END aoi222d4

MACRO aoi222d2
    CLASS CORE ;
    FOREIGN aoi222d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.370 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.910 0.800 2.310 ;
        RECT  0.120 1.460 0.500 2.310 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.670 2.000 2.070 ;
        RECT  1.180 1.460 1.620 2.070 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.700 2.840 2.100 ;
        RECT  2.300 1.700 2.740 2.460 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.506  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.020 4.040 2.630 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.527  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.340 2.020 4.980 2.630 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.618  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.710 3.700 6.660 4.140 ;
        RECT  5.710 3.340 6.360 4.140 ;
        RECT  5.710 1.700 5.950 4.140 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  6.700 4.450 7.100 5.600 ;
        RECT  5.390 4.450 5.790 5.600 ;
        RECT  4.030 4.340 4.430 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.370 0.000 6.770 0.980 ;
        RECT  4.780 0.000 5.180 0.980 ;
        RECT  2.690 0.000 3.090 0.980 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 4.260 3.130 4.500 ;
        RECT  1.990 3.300 4.990 3.540 ;
        RECT  1.350 0.980 2.450 1.220 ;
        RECT  2.210 1.220 6.430 1.460 ;
        RECT  6.190 1.220 6.430 2.550 ;
        RECT  6.190 2.310 7.240 2.550 ;
        RECT  0.720 3.260 1.120 4.020 ;
        RECT  5.230 1.220 5.470 4.020 ;
        RECT  0.720 3.780 5.470 4.020 ;
        RECT  7.110 1.000 7.510 1.940 ;
        RECT  6.190 2.860 7.720 3.100 ;
        RECT  7.480 1.630 7.720 3.710 ;
        RECT  7.270 2.860 7.720 3.710 ;
    END
END aoi222d2

MACRO aoi222d1
    CLASS CORE ;
    FOREIGN aoi222d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.520 0.550 2.920 ;
        RECT  0.120 2.520 0.500 3.580 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.460 1.460 2.180 1.900 ;
        RECT  1.300 2.140 1.700 2.540 ;
        RECT  1.460 1.460 1.700 2.540 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.980 2.580 2.740 3.020 ;
        RECT  1.980 2.140 2.380 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.502  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.980 2.700 3.860 3.100 ;
        RECT  3.420 2.580 3.860 3.100 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.532  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.540 2.020 4.980 2.460 ;
        RECT  3.220 2.020 4.980 2.340 ;
        RECT  3.220 1.940 3.620 2.340 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.515  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.100 2.700 5.480 3.580 ;
        RECT  4.630 2.700 5.480 3.100 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.073  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.240 4.570 1.480 ;
        RECT  2.490 0.980 2.730 1.480 ;
        RECT  0.930 0.980 2.730 1.220 ;
        RECT  0.620 1.460 1.170 1.900 ;
        RECT  0.930 0.980 1.170 1.900 ;
        RECT  0.750 3.260 1.150 3.660 ;
        RECT  0.790 1.460 1.060 3.660 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.970 4.440 5.370 5.600 ;
        RECT  3.550 4.440 3.950 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  2.970 0.000 3.370 0.980 ;
        RECT  0.290 0.000 0.690 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 4.130 3.200 4.370 ;
        RECT  2.230 3.440 4.520 3.680 ;
    END
END aoi222d1

MACRO aoi2222d4
    CLASS CORE ;
    FOREIGN aoi2222d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.385  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.370 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.406  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.840 0.860 2.240 ;
        RECT  0.120 1.460 0.500 2.240 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.529  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.710 2.580 2.180 3.020 ;
        RECT  1.710 2.040 2.110 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.580 2.580 3.300 3.020 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.960 1.460 10.580 1.900 ;
        RECT  9.810 2.540 10.210 2.940 ;
        RECT  9.960 1.460 10.210 2.940 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.700 2.140 11.080 3.580 ;
        RECT  10.550 2.140 11.080 2.540 ;
        END
    END C2
    PIN D1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 1.940 9.470 2.460 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 2.060 8.300 2.460 ;
        RECT  7.340 2.020 7.780 2.460 ;
        END
    END D2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.754  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.040 1.710 5.960 2.110 ;
        RECT  4.040 3.050 5.740 3.580 ;
        RECT  4.040 1.710 4.280 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  8.750 4.340 9.150 5.600 ;
        RECT  7.270 3.940 7.670 5.600 ;
        RECT  5.900 4.530 6.300 5.600 ;
        RECT  4.600 4.530 5.000 5.600 ;
        RECT  3.300 4.530 3.700 5.600 ;
        RECT  2.030 4.450 2.430 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  10.630 0.000 11.030 1.220 ;
        RECT  8.120 0.000 8.520 1.220 ;
        RECT  6.140 0.000 6.540 1.420 ;
        RECT  4.840 0.000 5.240 1.400 ;
        RECT  3.540 0.000 3.940 1.400 ;
        RECT  2.640 0.000 3.040 1.220 ;
        RECT  0.210 0.000 0.610 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.460 3.760 3.170 4.000 ;
        RECT  1.460 3.760 1.860 4.160 ;
        RECT  0.150 4.090 1.690 4.330 ;
        RECT  0.150 4.090 0.550 4.620 ;
        RECT  1.440 1.400 1.840 1.800 ;
        RECT  1.440 1.480 3.200 1.800 ;
        RECT  2.960 1.480 3.200 2.330 ;
        RECT  2.960 1.930 3.780 2.330 ;
        RECT  3.540 1.930 3.780 3.520 ;
        RECT  0.720 3.280 3.780 3.520 ;
        RECT  0.720 3.280 1.120 3.850 ;
        RECT  6.780 1.020 7.820 1.420 ;
        RECT  5.110 2.370 7.020 2.770 ;
        RECT  6.780 1.020 7.020 3.670 ;
        RECT  6.680 3.270 7.080 3.670 ;
        RECT  9.320 1.210 9.720 1.700 ;
        RECT  8.540 1.460 9.720 1.700 ;
        RECT  7.320 2.740 8.780 3.140 ;
        RECT  8.540 1.460 8.780 3.420 ;
        RECT  8.540 3.180 10.460 3.420 ;
        RECT  10.060 3.180 10.460 3.820 ;
        RECT  8.010 3.660 9.720 4.060 ;
        RECT  9.390 3.660 9.720 4.490 ;
        RECT  9.390 4.090 11.030 4.490 ;
        RECT  8.010 3.660 8.410 4.620 ;
    END
END aoi2222d4

MACRO aoi2222d2
    CLASS CORE ;
    FOREIGN aoi2222d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.385  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.370 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.406  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.840 0.860 2.240 ;
        RECT  0.120 1.460 0.500 2.240 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.529  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.710 2.580 2.180 3.020 ;
        RECT  1.710 2.040 2.110 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.900 2.580 3.300 3.200 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.790 1.460 9.460 1.900 ;
        RECT  8.640 2.540 9.040 2.940 ;
        RECT  8.790 1.460 9.040 2.940 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.580 2.140 9.960 3.580 ;
        RECT  9.380 2.140 9.960 2.540 ;
        END
    END C2
    PIN D1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.900 1.940 8.340 2.540 ;
        END
    END D1
    PIN D2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.220 2.020 7.180 2.460 ;
        END
    END D2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.482  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.100 3.050 4.980 3.580 ;
        RECT  4.100 1.710 4.790 2.110 ;
        RECT  4.100 1.710 4.340 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.080 5.600 ;
        RECT  7.580 4.340 7.980 5.600 ;
        RECT  6.100 3.940 6.500 5.600 ;
        RECT  4.730 4.530 5.130 5.600 ;
        RECT  3.430 4.530 3.830 5.600 ;
        RECT  2.030 4.450 2.430 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.080 0.740 ;
        RECT  9.460 0.000 9.860 1.220 ;
        RECT  6.950 0.000 7.350 1.220 ;
        RECT  4.970 0.000 5.370 1.420 ;
        RECT  3.490 0.000 3.890 1.420 ;
        RECT  2.640 0.000 3.040 1.220 ;
        RECT  0.210 0.000 0.610 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.460 3.760 3.170 4.160 ;
        RECT  0.150 4.090 1.690 4.330 ;
        RECT  0.150 4.090 0.550 4.620 ;
        RECT  1.440 1.400 1.840 1.800 ;
        RECT  1.440 1.480 2.660 1.800 ;
        RECT  2.420 1.930 3.300 2.330 ;
        RECT  2.420 1.480 2.660 3.520 ;
        RECT  0.720 3.280 2.660 3.520 ;
        RECT  0.720 3.280 1.120 3.850 ;
        RECT  5.610 1.020 6.650 1.420 ;
        RECT  4.580 2.370 5.850 2.770 ;
        RECT  5.610 1.020 5.850 3.670 ;
        RECT  5.510 3.270 5.910 3.670 ;
        RECT  8.150 1.210 8.550 1.700 ;
        RECT  7.420 1.460 8.550 1.700 ;
        RECT  6.150 2.740 7.660 3.140 ;
        RECT  7.420 1.460 7.660 3.420 ;
        RECT  7.420 3.180 9.290 3.420 ;
        RECT  8.890 3.180 9.290 3.820 ;
        RECT  6.840 3.660 8.550 4.060 ;
        RECT  8.220 3.660 8.550 4.490 ;
        RECT  8.220 4.090 9.860 4.490 ;
        RECT  6.840 3.660 7.240 4.620 ;
    END
END aoi2222d2

MACRO aoi2222d1
    CLASS CORE ;
    FOREIGN aoi2222d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.340 1.940 7.780 2.540 ;
        END
    END D1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.385  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.370 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.406  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.840 0.860 2.240 ;
        RECT  0.120 1.460 0.500 2.240 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.529  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.710 2.580 2.180 3.020 ;
        RECT  1.710 2.040 2.110 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.900 2.580 3.300 3.200 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.230 1.460 8.900 1.900 ;
        RECT  8.080 2.540 8.480 2.940 ;
        RECT  8.230 1.460 8.480 2.940 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.391  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 2.140 9.400 3.580 ;
        RECT  8.820 2.140 9.400 2.540 ;
        END
    END C2
    PIN D2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 2.060 6.570 2.460 ;
        RECT  5.660 2.020 6.100 2.460 ;
        END
    END D2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.540 3.050 4.420 3.580 ;
        RECT  3.540 1.710 4.230 2.110 ;
        RECT  3.540 1.710 3.780 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 9.520 5.600 ;
        RECT  7.020 4.340 7.420 5.600 ;
        RECT  5.540 3.940 5.940 5.600 ;
        RECT  4.170 4.530 4.570 5.600 ;
        RECT  2.030 4.450 2.430 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 9.520 0.740 ;
        RECT  8.900 0.000 9.300 1.220 ;
        RECT  6.390 0.000 6.790 1.220 ;
        RECT  4.410 0.000 4.810 1.420 ;
        RECT  2.640 0.000 3.040 1.220 ;
        RECT  0.210 0.000 0.610 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.460 3.760 3.170 4.160 ;
        RECT  0.150 4.090 1.690 4.330 ;
        RECT  0.150 4.090 0.550 4.620 ;
        RECT  1.440 1.400 1.840 1.800 ;
        RECT  1.440 1.480 2.660 1.800 ;
        RECT  2.420 1.930 3.300 2.330 ;
        RECT  2.420 1.480 2.660 3.520 ;
        RECT  0.720 3.280 2.660 3.520 ;
        RECT  0.720 3.280 1.120 3.850 ;
        RECT  5.050 1.020 6.090 1.420 ;
        RECT  4.020 2.370 5.290 2.770 ;
        RECT  5.050 1.020 5.290 3.670 ;
        RECT  4.950 3.270 5.350 3.670 ;
        RECT  7.590 1.210 7.990 1.700 ;
        RECT  6.810 1.460 7.990 1.700 ;
        RECT  5.590 2.740 7.050 3.140 ;
        RECT  6.810 1.460 7.050 3.420 ;
        RECT  6.810 3.180 8.730 3.420 ;
        RECT  8.330 3.180 8.730 3.820 ;
        RECT  6.280 3.660 7.990 4.060 ;
        RECT  7.660 3.660 7.990 4.490 ;
        RECT  7.660 4.090 9.300 4.490 ;
        RECT  6.280 3.660 6.680 4.620 ;
    END
END aoi2222d1

MACRO aoi221d4
    CLASS CORE ;
    FOREIGN aoi221d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.503  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.860 1.080 2.460 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.320 2.580 2.180 2.940 ;
        RECT  1.320 2.520 1.720 2.940 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.940 3.300 2.460 ;
        RECT  2.240 1.940 3.300 2.340 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.493  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.220 3.480 3.580 ;
        RECT  3.080 2.700 3.480 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.780 2.020 4.420 2.460 ;
        RECT  3.780 2.020 4.180 3.270 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.942  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.510 3.270 6.910 4.570 ;
        RECT  4.920 1.700 6.830 1.940 ;
        RECT  4.920 3.270 6.910 3.580 ;
        RECT  4.920 3.140 5.730 3.580 ;
        RECT  4.920 1.700 5.160 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  7.250 4.380 7.650 5.600 ;
        RECT  4.560 4.500 4.960 5.600 ;
        RECT  3.290 4.620 3.690 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.170 0.000 7.570 0.980 ;
        RECT  5.860 0.000 6.260 0.980 ;
        RECT  4.510 0.000 4.910 0.980 ;
        RECT  2.010 0.000 2.410 0.980 ;
        RECT  0.150 0.000 0.550 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 4.100 1.120 4.620 ;
        RECT  0.720 4.380 2.390 4.620 ;
        RECT  1.420 3.490 1.820 4.060 ;
        RECT  1.420 3.820 4.430 4.060 ;
        RECT  2.730 3.820 4.430 4.220 ;
        RECT  0.770 1.220 7.370 1.460 ;
        RECT  0.120 1.380 1.170 1.620 ;
        RECT  7.130 1.220 7.370 2.550 ;
        RECT  7.130 2.150 7.760 2.550 ;
        RECT  0.120 1.380 0.360 3.450 ;
        RECT  0.120 3.050 0.550 3.450 ;
        RECT  7.850 1.510 8.250 1.910 ;
        RECT  5.950 2.520 6.890 3.030 ;
        RECT  5.950 2.790 8.250 3.030 ;
        RECT  8.000 1.510 8.250 3.450 ;
        RECT  7.820 2.790 8.250 3.450 ;
    END
END aoi221d4

MACRO aoi221d2
    CLASS CORE ;
    FOREIGN aoi221d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.509  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.020 1.080 2.810 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.320 2.580 2.180 3.020 ;
        RECT  1.320 2.520 1.720 3.020 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.470  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.960 3.300 2.460 ;
        RECT  2.290 1.960 3.300 2.360 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.190 3.140 3.860 3.580 ;
        RECT  3.190 2.700 3.590 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.490  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.070 2.020 4.470 3.020 ;
        RECT  3.980 2.020 4.470 2.460 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.671  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 3.350 6.100 4.140 ;
        RECT  5.030 3.350 6.100 3.750 ;
        RECT  5.030 1.700 5.590 2.100 ;
        RECT  5.030 1.700 5.270 3.750 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.150 4.450 6.550 5.600 ;
        RECT  4.840 4.450 5.240 5.600 ;
        RECT  3.490 4.620 3.890 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  6.050 0.000 6.450 0.980 ;
        RECT  4.590 0.000 4.990 0.980 ;
        RECT  2.180 0.000 2.420 1.190 ;
        RECT  0.230 0.000 0.470 1.190 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.770 4.180 2.440 4.420 ;
        RECT  1.470 3.350 2.920 3.750 ;
        RECT  2.680 3.350 2.920 4.220 ;
        RECT  2.680 3.820 4.540 4.220 ;
        RECT  2.840 1.220 6.490 1.460 ;
        RECT  0.770 1.430 3.080 1.670 ;
        RECT  0.120 1.540 1.170 1.780 ;
        RECT  6.250 1.220 6.490 2.630 ;
        RECT  6.250 2.230 6.680 2.630 ;
        RECT  0.120 1.540 0.360 3.450 ;
        RECT  0.120 3.050 0.600 3.450 ;
        RECT  6.730 1.590 7.160 1.990 ;
        RECT  5.510 2.620 5.910 3.110 ;
        RECT  5.510 2.870 7.160 3.110 ;
        RECT  6.920 1.590 7.160 3.550 ;
        RECT  6.730 2.870 7.160 3.550 ;
    END
END aoi221d2

MACRO aoi221d1
    CLASS CORE ;
    FOREIGN aoi221d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.090 1.060 2.530 ;
        RECT  0.620 2.020 1.060 2.530 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.580 2.130 3.020 ;
        RECT  1.740 2.130 1.980 3.020 ;
        RECT  1.560 2.130 1.980 2.530 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.458  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.350 1.850 2.810 2.260 ;
        RECT  2.350 1.850 2.720 2.460 ;
        END
    END B2
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.580 3.860 3.020 ;
        RECT  2.980 2.580 3.860 2.920 ;
        RECT  2.980 2.520 3.380 2.920 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.476  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.940 4.360 2.340 ;
        RECT  3.980 1.460 4.360 2.340 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.608  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.320 0.980 4.330 1.220 ;
        RECT  1.310 1.220 3.560 1.460 ;
        RECT  0.120 1.540 1.710 1.780 ;
        RECT  1.310 1.220 1.710 1.780 ;
        RECT  0.120 3.140 0.500 4.040 ;
        RECT  0.120 1.540 0.360 4.040 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.360 4.180 3.760 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  2.680 0.000 3.080 0.980 ;
        RECT  0.340 0.000 0.740 1.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.050 4.160 2.450 4.610 ;
        RECT  0.760 4.370 2.450 4.610 ;
        RECT  1.260 2.940 1.500 3.870 ;
        RECT  1.260 3.470 4.330 3.870 ;
    END
END aoi221d1

MACRO aoi21d4
    CLASS CORE ;
    FOREIGN aoi21d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.920 0.980 2.740 1.260 ;
        RECT  1.840 1.890 2.160 2.290 ;
        RECT  1.920 0.980 2.160 2.290 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.416  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.710 3.010 1.500 3.250 ;
        RECT  0.710 2.320 1.010 3.250 ;
        RECT  0.700 1.460 1.000 2.620 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.457  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.900 0.470 3.300 ;
        RECT  0.120 2.020 0.460 3.300 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.957  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.680 3.050 5.450 3.580 ;
        RECT  3.740 1.770 5.450 2.170 ;
        RECT  4.660 1.770 4.900 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.470 4.260 4.880 5.600 ;
        RECT  3.180 4.300 3.580 5.600 ;
        RECT  0.740 4.180 1.140 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.480 0.000 4.880 1.150 ;
        RECT  3.180 0.000 3.580 1.120 ;
        RECT  0.150 0.000 0.550 1.270 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.170 3.570 1.720 3.810 ;
        RECT  1.480 3.570 1.720 4.620 ;
        RECT  1.480 4.220 1.950 4.620 ;
        RECT  1.430 1.020 1.670 1.720 ;
        RECT  1.330 1.500 1.570 2.770 ;
        RECT  1.330 2.530 2.960 2.770 ;
        RECT  2.560 2.410 2.960 2.810 ;
        RECT  1.960 2.530 2.200 3.980 ;
        RECT  1.960 3.740 2.690 3.980 ;
        RECT  2.290 3.740 2.690 4.620 ;
        RECT  2.400 1.770 3.440 2.170 ;
        RECT  3.200 2.410 3.890 2.810 ;
        RECT  3.200 1.770 3.440 3.450 ;
        RECT  2.440 3.050 3.440 3.450 ;
    END
END aoi21d4

MACRO aoi21d2
    CLASS CORE ;
    FOREIGN aoi21d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.425  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.050 2.020 2.740 2.460 ;
        RECT  2.050 1.730 2.450 2.460 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.900 1.330 2.300 ;
        RECT  0.120 1.460 0.500 2.300 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.580 1.060 3.050 ;
        RECT  0.400 2.580 1.060 2.980 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.593  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.360 3.140 4.980 3.580 ;
        RECT  4.540 1.460 4.980 3.580 ;
        RECT  4.310 1.460 4.980 1.860 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.980 4.710 5.380 5.600 ;
        RECT  3.620 4.710 4.020 5.600 ;
        RECT  0.790 4.710 1.190 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  5.050 0.000 5.450 1.160 ;
        RECT  3.660 0.000 4.060 1.160 ;
        RECT  1.990 0.000 2.390 0.900 ;
        RECT  0.150 0.000 0.550 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 3.290 1.850 3.530 ;
        RECT  1.400 1.190 1.810 1.590 ;
        RECT  1.570 1.190 1.810 2.940 ;
        RECT  2.980 2.540 3.380 2.940 ;
        RECT  1.570 2.700 3.380 2.940 ;
        RECT  2.240 2.700 2.640 3.540 ;
        RECT  2.890 1.380 3.290 1.780 ;
        RECT  2.890 1.540 4.020 1.780 ;
        RECT  3.780 2.100 4.300 2.500 ;
        RECT  3.780 1.540 4.020 3.580 ;
        RECT  2.940 3.180 4.020 3.580 ;
    END
END aoi21d2

MACRO aoi21d1
    CLASS CORE ;
    FOREIGN aoi21d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.230 1.060 3.020 ;
        END
    END A
    PIN B1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.419  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.460 2.180 1.900 ;
        RECT  1.420 2.230 1.850 2.630 ;
        RECT  1.610 1.460 1.850 2.630 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.120 2.580 2.680 3.020 ;
        RECT  2.120 2.180 2.520 3.020 ;
        END
    END B2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.146  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.590 1.370 1.990 ;
        RECT  0.120 3.340 0.610 4.140 ;
        RECT  0.120 1.590 0.360 4.140 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  1.620 4.100 2.020 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  2.200 0.000 2.600 1.220 ;
        RECT  0.320 0.000 0.720 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.950 3.530 2.650 3.770 ;
    END
END aoi21d1

MACRO aoi211d4
    CLASS CORE ;
    FOREIGN aoi211d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.494  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.500 2.180 2.940 2.580 ;
        RECT  2.360 3.140 2.740 3.580 ;
        RECT  2.500 2.180 2.740 3.580 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.800 2.180 2.260 2.580 ;
        RECT  1.800 2.180 2.150 3.020 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.120 2.510 1.560 2.910 ;
        RECT  1.180 2.020 1.560 2.910 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.421  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.900 0.820 3.300 ;
        RECT  0.120 2.020 0.500 3.300 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.964  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.800 3.050 6.570 3.580 ;
        RECT  4.860 1.730 6.570 2.130 ;
        RECT  5.310 1.730 5.550 3.580 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.590 4.260 6.000 5.600 ;
        RECT  4.300 4.300 4.700 5.600 ;
        RECT  0.790 4.100 1.190 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.600 0.000 6.000 1.150 ;
        RECT  4.300 0.000 4.700 1.430 ;
        RECT  2.150 0.000 2.550 1.300 ;
        RECT  0.170 0.000 0.570 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.170 3.540 1.870 3.780 ;
        RECT  1.370 1.380 1.770 1.780 ;
        RECT  1.370 1.540 3.190 1.780 ;
        RECT  2.790 1.650 3.420 1.940 ;
        RECT  3.180 2.400 3.640 2.790 ;
        RECT  3.180 1.650 3.420 3.300 ;
        RECT  2.980 3.040 3.220 4.500 ;
        RECT  2.790 4.100 3.220 4.500 ;
        RECT  3.560 1.040 3.960 1.440 ;
        RECT  3.720 1.040 3.960 2.100 ;
        RECT  3.880 2.390 5.010 2.790 ;
        RECT  3.880 1.800 4.120 4.140 ;
        RECT  3.560 3.740 4.120 4.140 ;
    END
END aoi211d4

MACRO aoi211d2
    CLASS CORE ;
    FOREIGN aoi211d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.443  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 2.180 3.300 3.020 ;
        RECT  2.590 2.180 3.300 2.580 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.480  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.110 3.220 2.740 3.500 ;
        RECT  2.110 2.520 2.350 3.500 ;
        RECT  1.860 2.520 2.350 2.920 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.580 1.620 3.020 ;
        RECT  0.980 2.500 1.380 2.900 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.180 0.550 2.580 ;
        RECT  0.120 2.180 0.500 3.020 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.417  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.890 3.110 5.540 3.580 ;
        RECT  4.890 3.050 5.410 3.580 ;
        RECT  5.170 1.380 5.410 3.580 ;
        RECT  4.870 1.380 5.410 1.780 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.500 4.260 5.910 5.600 ;
        RECT  4.120 4.710 4.520 5.600 ;
        RECT  0.790 4.100 1.190 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  5.610 0.000 6.010 1.150 ;
        RECT  4.250 0.000 4.650 0.890 ;
        RECT  2.010 0.000 2.410 1.300 ;
        RECT  0.170 0.000 0.570 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.170 3.540 1.870 3.780 ;
        RECT  1.420 1.700 3.930 1.940 ;
        RECT  3.690 1.700 3.930 3.500 ;
        RECT  2.980 3.260 3.930 3.500 ;
        RECT  2.980 3.260 3.220 4.150 ;
        RECT  2.830 3.750 3.220 4.150 ;
        RECT  3.480 1.160 4.410 1.400 ;
        RECT  4.170 2.030 4.930 2.430 ;
        RECT  4.170 1.160 4.410 4.060 ;
        RECT  3.530 3.820 4.410 4.060 ;
    END
END aoi211d2

MACRO aoi211d1
    CLASS CORE ;
    FOREIGN aoi211d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.462  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.020 1.060 2.810 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.497  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.300 2.500 1.700 2.900 ;
        RECT  1.180 3.110 1.620 3.580 ;
        RECT  1.300 2.500 1.620 3.580 ;
        END
    END B
    PIN C1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.880 3.180 2.740 3.580 ;
        RECT  2.300 3.140 2.740 3.580 ;
        END
    END C1
    PIN C2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.560 2.500 3.240 2.900 ;
        RECT  2.860 2.020 3.240 2.900 ;
        END
    END C2
    PIN ZN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.593  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.540 1.130 2.180 2.050 ;
        RECT  0.120 1.130 2.180 1.370 ;
        RECT  0.120 3.050 0.550 3.450 ;
        RECT  0.120 1.080 0.550 1.500 ;
        RECT  0.120 1.080 0.360 3.450 ;
        END
    END ZN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.160 4.380 2.560 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.810 0.000 3.210 1.430 ;
        RECT  0.920 0.000 1.320 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.360 3.850 3.210 4.090 ;
        RECT  1.360 3.850 1.760 4.500 ;
    END
END aoi211d1

MACRO an12d4
    CLASS CORE ;
    FOREIGN an12d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.990 0.540 3.400 ;
        RECT  0.130 2.550 0.500 3.400 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.130 2.370 3.580 ;
        RECT  2.130 2.520 2.370 3.580 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.100  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.100 3.130 4.810 3.370 ;
        RECT  3.100 1.630 4.810 1.870 ;
        RECT  3.980 3.130 4.420 3.580 ;
        RECT  4.180 1.630 4.420 3.580 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.840 4.620 4.240 5.600 ;
        RECT  2.470 4.620 2.870 5.600 ;
        RECT  1.000 4.340 1.240 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.840 0.000 4.240 0.980 ;
        RECT  2.470 0.000 2.870 0.890 ;
        RECT  0.540 0.000 0.780 1.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.460 1.820 1.140 2.060 ;
        RECT  0.900 1.820 1.140 3.890 ;
        RECT  0.150 3.650 1.140 3.890 ;
        RECT  1.240 1.340 2.850 1.580 ;
        RECT  2.610 2.510 3.940 2.810 ;
        RECT  2.610 1.340 2.850 4.090 ;
        RECT  1.690 3.850 2.850 4.090 ;
    END
END an12d4

MACRO an12d2
    CLASS CORE ;
    FOREIGN an12d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.990 0.540 3.400 ;
        RECT  0.130 2.550 0.500 3.400 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.990 2.350 3.580 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.272  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.100 3.530 3.860 3.930 ;
        RECT  3.620 1.370 3.860 3.930 ;
        RECT  3.400 3.130 3.860 3.930 ;
        RECT  3.100 1.370 3.860 1.610 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.840 4.620 4.240 5.600 ;
        RECT  2.470 4.620 2.870 5.600 ;
        RECT  1.000 4.330 1.240 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  3.840 0.000 4.240 0.980 ;
        RECT  2.470 0.000 2.870 0.890 ;
        RECT  0.540 0.000 0.780 1.430 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.460 1.850 1.140 2.090 ;
        RECT  0.900 1.850 1.140 3.890 ;
        RECT  0.150 3.650 1.140 3.890 ;
        RECT  1.240 1.050 1.620 1.450 ;
        RECT  1.380 1.050 1.620 2.750 ;
        RECT  1.380 2.510 3.250 2.750 ;
        RECT  2.590 2.510 3.250 2.780 ;
        RECT  2.590 2.510 2.830 4.090 ;
        RECT  1.690 3.850 2.830 4.090 ;
    END
END an12d2

MACRO an12d1
    CLASS CORE ;
    FOREIGN an12d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.990 0.540 3.400 ;
        RECT  0.130 2.550 0.500 3.400 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.580 3.580 ;
        RECT  2.160 2.990 2.580 3.580 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.087  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.410 1.290 3.800 3.930 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  2.700 4.620 3.100 5.600 ;
        RECT  1.230 4.330 1.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  2.710 0.000 3.110 0.890 ;
        RECT  0.540 0.000 0.780 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.460 1.840 1.500 2.080 ;
        RECT  1.260 1.840 1.500 3.890 ;
        RECT  0.380 3.650 1.500 3.890 ;
        RECT  1.240 1.130 3.160 1.370 ;
        RECT  2.920 1.130 3.160 4.090 ;
        RECT  1.920 3.850 3.160 4.090 ;
    END
END an12d1

MACRO an04da
    CLASS CORE ;
    FOREIGN an04da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.410 0.810 2.650 ;
        RECT  0.120 1.740 0.500 2.650 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.320 3.040 1.500 3.580 ;
        RECT  1.080 2.960 1.500 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.500 2.180 2.840 ;
        RECT  1.180 2.500 2.180 2.730 ;
        RECT  1.180 2.020 1.620 2.730 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.810 3.580 ;
        RECT  2.570 2.820 2.810 3.580 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.760  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.850 1.130 8.280 3.450 ;
        RECT  4.790 1.130 8.280 3.310 ;
        RECT  4.790 1.130 6.410 4.300 ;
        RECT  3.670 2.540 8.280 3.070 ;
        RECT  4.550 1.130 8.280 3.070 ;
        RECT  3.230 1.130 8.280 1.630 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.400 5.600 ;
        RECT  6.750 3.540 7.150 5.600 ;
        RECT  5.260 4.620 5.670 5.600 ;
        RECT  4.150 3.300 4.550 5.600 ;
        RECT  2.810 4.620 3.210 5.600 ;
        RECT  1.460 4.620 1.860 5.600 ;
        RECT  0.150 4.020 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.400 0.740 ;
        RECT  7.080 0.000 7.480 0.890 ;
        RECT  5.540 0.000 5.940 0.890 ;
        RECT  4.000 0.000 4.400 0.890 ;
        RECT  2.490 0.000 2.890 1.520 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 0.970 2.260 1.510 ;
        RECT  1.860 0.970 2.260 2.270 ;
        RECT  1.860 1.860 4.320 2.270 ;
        RECT  2.980 1.860 4.320 2.310 ;
        RECT  3.040 1.860 3.440 4.310 ;
        RECT  0.900 3.810 3.440 4.310 ;
    END
END an04da

MACRO an04d7
    CLASS CORE ;
    FOREIGN an04d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.486  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.410 0.810 2.650 ;
        RECT  0.120 1.740 0.500 2.650 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.486  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.040 1.500 3.580 ;
        RECT  1.080 2.810 1.500 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.477  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.280 2.170 2.520 ;
        RECT  1.180 2.020 1.620 2.520 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.486  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.770 3.580 ;
        RECT  2.530 2.820 2.770 3.580 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.732  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.550 2.450 7.160 2.850 ;
        RECT  6.780 1.130 7.160 2.850 ;
        RECT  3.650 1.130 7.160 1.530 ;
        RECT  6.160 2.450 6.560 3.450 ;
        RECT  4.750 2.450 4.990 4.210 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.730 3.730 7.130 5.600 ;
        RECT  5.420 3.690 5.820 5.600 ;
        RECT  3.940 3.210 4.510 3.450 ;
        RECT  3.940 3.210 4.180 5.600 ;
        RECT  2.770 4.620 3.170 5.600 ;
        RECT  1.460 4.560 1.860 5.600 ;
        RECT  0.150 3.950 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  5.960 0.000 6.360 0.890 ;
        RECT  4.420 0.000 4.820 0.890 ;
        RECT  2.690 0.000 3.090 1.520 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.120 2.100 1.360 ;
        RECT  1.860 1.120 2.100 2.040 ;
        RECT  1.860 1.760 3.260 2.040 ;
        RECT  3.020 1.790 6.400 2.190 ;
        RECT  0.900 3.950 1.460 4.190 ;
        RECT  3.020 1.760 3.260 4.260 ;
        RECT  1.220 4.020 3.260 4.260 ;
    END
END an04d7

MACRO an04d4
    CLASS CORE ;
    FOREIGN an04d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.490 0.670 2.900 ;
        RECT  0.120 2.020 0.490 2.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 3.140 1.620 3.580 ;
        RECT  1.220 2.530 1.460 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.960 2.020 2.200 2.870 ;
        RECT  1.740 2.020 2.200 2.460 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.140 2.980 3.580 ;
        RECT  2.740 2.530 2.980 3.580 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.718  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.730 3.140 5.450 3.380 ;
        RECT  3.740 1.730 5.450 1.970 ;
        RECT  4.540 1.730 4.980 3.380 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.600 5.600 ;
        RECT  4.560 4.320 4.800 5.600 ;
        RECT  3.260 4.320 3.500 5.600 ;
        RECT  1.640 4.710 2.040 5.600 ;
        RECT  0.230 4.040 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.600 0.740 ;
        RECT  4.390 0.000 4.630 1.130 ;
        RECT  3.080 0.000 3.320 1.130 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 1.540 3.490 1.780 ;
        RECT  3.250 2.510 4.070 2.750 ;
        RECT  3.250 1.540 3.490 4.060 ;
        RECT  0.890 3.820 3.490 4.060 ;
    END
END an04d4

MACRO an04d2
    CLASS CORE ;
    FOREIGN an04d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.490 0.670 2.900 ;
        RECT  0.120 2.020 0.490 2.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.330 3.580 ;
        RECT  1.090 2.740 1.330 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.020 2.010 3.160 ;
        RECT  1.180 2.020 2.010 2.460 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.180 2.740 3.020 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.266  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  3.580 1.060 3.820 4.140 ;
        RECT  3.370 1.060 3.820 1.460 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  4.330 3.900 4.570 5.600 ;
        RECT  2.910 4.710 3.310 5.600 ;
        RECT  1.430 4.480 1.670 5.600 ;
        RECT  0.250 4.480 0.490 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  4.200 0.000 4.440 1.470 ;
        RECT  2.680 0.000 2.920 1.230 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 1.540 2.540 1.780 ;
        RECT  2.300 1.700 3.320 1.940 ;
        RECT  3.080 1.700 3.320 3.450 ;
        RECT  2.940 3.210 3.180 4.060 ;
        RECT  0.760 3.820 3.180 4.060 ;
    END
END an04d2

MACRO an04d1
    CLASS CORE ;
    FOREIGN an04d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.490 0.670 2.900 ;
        RECT  0.120 2.020 0.490 2.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.330 3.580 ;
        RECT  1.090 2.740 1.330 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.020 2.010 3.160 ;
        RECT  1.180 2.020 2.010 2.460 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.180 2.740 3.020 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.177  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.860 4.140 ;
        RECT  3.620 1.060 3.860 4.140 ;
        RECT  3.440 1.060 3.860 1.460 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  2.910 4.710 3.310 5.600 ;
        RECT  1.430 4.480 1.670 5.600 ;
        RECT  0.250 4.480 0.490 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  2.680 0.000 2.920 1.230 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 1.540 2.540 1.780 ;
        RECT  2.300 1.700 3.320 1.940 ;
        RECT  3.080 1.700 3.320 3.450 ;
        RECT  2.940 3.210 3.180 4.060 ;
        RECT  0.760 3.820 3.180 4.060 ;
    END
END an04d1

MACRO an04d0
    CLASS CORE ;
    FOREIGN an04d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.490 0.840 2.900 ;
        RECT  0.120 2.020 0.490 2.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.460 3.380 ;
        RECT  1.220 2.740 1.460 3.380 ;
        RECT  0.620 3.140 1.060 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.140 2.180 3.580 ;
        RECT  1.900 2.730 2.180 3.580 ;
        END
    END A3
    PIN A4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.500 2.020 2.900 2.580 ;
        RECT  2.300 2.020 2.900 2.500 ;
        END
    END A4
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.669  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 3.700 3.990 4.140 ;
        RECT  3.740 1.610 3.990 4.140 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 4.480 5.600 ;
        RECT  3.100 4.380 3.340 5.600 ;
        RECT  1.430 4.480 1.670 5.600 ;
        RECT  0.250 4.480 0.490 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 4.480 0.740 ;
        RECT  2.880 0.000 3.120 1.230 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 1.540 3.500 1.780 ;
        RECT  3.260 1.540 3.500 3.450 ;
        RECT  2.940 3.210 3.500 3.450 ;
        RECT  2.940 3.210 3.180 4.060 ;
        RECT  0.760 3.820 3.180 4.060 ;
    END
END an04d0

MACRO an03da
    CLASS CORE ;
    FOREIGN an03da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.440 0.800 2.850 ;
        RECT  0.120 1.900 0.500 2.850 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.090 2.330 1.620 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.860 2.510 2.740 3.020 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.748  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.800 3.820 7.680 4.320 ;
        RECT  4.110 1.240 7.680 4.320 ;
        RECT  2.840 1.220 7.280 1.720 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  7.260 4.550 7.660 5.600 ;
        RECT  5.960 4.550 6.360 5.600 ;
        RECT  4.660 4.550 5.060 5.600 ;
        RECT  3.360 4.550 3.760 5.600 ;
        RECT  2.060 4.180 2.460 5.600 ;
        RECT  0.720 4.180 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  6.540 0.000 6.940 0.990 ;
        RECT  5.060 0.000 5.460 0.990 ;
        RECT  3.580 0.000 3.980 0.990 ;
        RECT  1.980 0.000 2.380 0.990 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.230 2.580 1.630 ;
        RECT  2.180 1.230 2.580 2.280 ;
        RECT  2.180 1.950 3.880 2.280 ;
        RECT  2.970 1.950 3.880 2.350 ;
        RECT  2.970 1.950 3.370 3.590 ;
        RECT  0.150 3.260 3.370 3.590 ;
        RECT  0.150 3.260 1.860 3.660 ;
        RECT  0.150 3.260 0.550 3.850 ;
        RECT  1.460 3.260 1.860 3.940 ;
    END
END an03da

MACRO an03d7
    CLASS CORE ;
    FOREIGN an03d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.470 0.800 2.880 ;
        RECT  0.120 1.820 0.500 2.880 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.477  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.070 2.520 1.620 3.020 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.860 2.410 2.740 3.020 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.942  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.780 1.230 6.140 1.470 ;
        RECT  2.780 3.880 5.780 4.120 ;
        RECT  5.100 2.580 5.540 3.020 ;
        RECT  5.190 1.230 5.430 4.120 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  6.160 3.730 6.560 5.600 ;
        RECT  4.640 4.550 5.040 5.600 ;
        RECT  3.340 4.550 3.740 5.600 ;
        RECT  2.020 4.310 2.420 5.600 ;
        RECT  0.800 4.110 1.040 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.000 0.000 5.400 0.990 ;
        RECT  3.520 0.000 3.920 0.990 ;
        RECT  2.030 0.000 2.270 1.420 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.230 1.790 1.470 ;
        RECT  1.550 1.230 1.790 2.120 ;
        RECT  1.550 1.720 4.950 2.120 ;
        RECT  3.240 1.720 3.480 3.500 ;
        RECT  0.150 3.260 3.480 3.500 ;
    END
END an03d7

MACRO an03d4
    CLASS CORE ;
    FOREIGN an03d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.460 2.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 1.620 2.460 ;
        RECT  1.180 2.020 1.500 2.890 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.481  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.050 2.320 3.590 ;
        RECT  1.990 2.520 2.320 3.590 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.760 4.810 3.450 ;
        RECT  3.260 2.580 4.810 3.020 ;
        RECT  3.260 1.760 3.500 3.450 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 5.040 5.600 ;
        RECT  3.900 4.620 4.300 5.600 ;
        RECT  2.590 4.620 2.990 5.600 ;
        RECT  1.000 4.270 1.240 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 5.040 0.740 ;
        RECT  3.750 0.000 4.160 1.020 ;
        RECT  2.410 0.000 2.820 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 2.100 1.780 ;
        RECT  1.860 1.540 2.100 2.280 ;
        RECT  1.860 2.040 3.020 2.280 ;
        RECT  2.780 2.040 3.020 2.890 ;
        RECT  0.700 1.540 0.940 4.030 ;
        RECT  0.150 3.790 1.600 4.030 ;
        RECT  1.380 3.830 2.140 4.070 ;
    END
END an03d4

MACRO an03d2
    CLASS CORE ;
    FOREIGN an03d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.540 2.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.780 2.700 1.480 2.940 ;
        RECT  0.620 3.140 1.060 3.580 ;
        RECT  0.780 2.700 1.060 3.580 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.930 2.000 2.460 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.203  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.800 3.140 3.300 3.780 ;
        RECT  2.880 1.390 3.120 3.780 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  3.440 4.300 3.690 5.600 ;
        RECT  2.110 4.480 2.350 5.600 ;
        RECT  1.180 4.680 1.580 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  3.370 0.000 3.780 1.020 ;
        RECT  1.960 0.000 2.370 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.210 2.620 1.450 ;
        RECT  2.380 1.210 2.620 2.940 ;
        RECT  2.050 2.700 2.620 2.940 ;
        RECT  1.180 3.790 2.290 4.030 ;
        RECT  2.050 2.700 2.290 4.030 ;
        RECT  0.710 3.860 1.420 4.100 ;
        RECT  0.710 3.860 0.950 4.570 ;
        RECT  0.150 4.330 0.950 4.570 ;
    END
END an03d2

MACRO an03d1
    CLASS CORE ;
    FOREIGN an03d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.020 0.540 2.900 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.490 3.500 ;
        RECT  1.080 2.820 1.490 3.500 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 2.000 2.460 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.034  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.390 3.240 3.780 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.290 4.480 2.530 5.600 ;
        RECT  1.180 4.630 1.580 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.060 0.000 2.460 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.210 2.620 1.450 ;
        RECT  2.380 1.210 2.620 4.030 ;
        RECT  0.150 3.790 2.620 4.030 ;
    END
END an03d1

MACRO an03d0
    CLASS CORE ;
    FOREIGN an03d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.930 0.540 2.910 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 3.140 1.480 3.500 ;
        RECT  1.080 2.810 1.480 3.500 ;
        END
    END A2
    PIN A3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.020 2.000 2.460 ;
        END
    END A3
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.936  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.400 3.240 4.620 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.180 4.480 2.420 5.600 ;
        RECT  1.180 4.660 1.580 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  1.960 0.000 2.360 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.210 2.640 1.450 ;
        RECT  2.400 1.210 2.640 4.030 ;
        RECT  0.150 3.790 2.640 4.030 ;
    END
END an03d0

MACRO an02da
    CLASS CORE ;
    FOREIGN an02da 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.485  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.080 0.800 2.600 ;
        RECT  0.120 2.020 0.500 2.460 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.477  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.080 1.850 1.540 2.460 ;
        RECT  1.080 1.850 1.480 2.700 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.510  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.580 7.160 3.020 ;
        RECT  6.730 1.170 7.130 1.570 ;
        RECT  6.160 1.210 6.970 3.290 ;
        RECT  6.160 1.210 6.560 3.450 ;
        RECT  3.500 1.210 6.970 3.030 ;
        RECT  4.940 1.210 5.440 4.340 ;
        RECT  3.640 1.210 4.070 4.580 ;
        RECT  2.340 2.540 4.070 3.040 ;
        RECT  2.380 1.210 6.970 1.680 ;
        RECT  2.340 2.540 2.770 4.050 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.280 5.600 ;
        RECT  6.730 3.740 7.130 5.600 ;
        RECT  5.420 4.620 5.820 5.600 ;
        RECT  4.300 3.260 4.700 5.600 ;
        RECT  3.000 3.500 3.400 5.600 ;
        RECT  1.490 4.150 1.890 5.600 ;
        RECT  0.150 3.050 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.280 0.740 ;
        RECT  5.990 0.000 6.390 0.980 ;
        RECT  4.590 0.000 4.990 0.980 ;
        RECT  3.120 0.000 3.520 0.980 ;
        RECT  1.780 0.000 2.180 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 1.110 1.470 1.620 ;
        RECT  0.230 1.120 2.100 1.620 ;
        RECT  1.770 1.120 2.100 3.440 ;
        RECT  1.770 1.910 3.270 2.310 ;
        RECT  1.770 1.910 2.110 3.440 ;
        RECT  0.820 2.940 2.110 3.440 ;
        RECT  0.820 2.940 1.260 4.100 ;
    END
END an02da

MACRO an02d7
    CLASS CORE ;
    FOREIGN an02d7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.532  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.320 0.800 2.720 ;
        RECT  0.120 2.020 0.500 2.720 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.060 2.020 1.620 2.510 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.206  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.310 1.210 5.980 1.450 ;
        RECT  3.420 2.050 5.550 2.290 ;
        RECT  5.310 1.210 5.550 2.290 ;
        RECT  5.070 2.050 5.310 4.130 ;
        RECT  4.170 0.980 4.410 2.290 ;
        RECT  3.750 2.050 3.990 3.870 ;
        RECT  2.630 2.930 3.990 3.170 ;
        RECT  3.420 2.020 3.860 3.170 ;
        RECT  3.240 1.370 3.480 2.270 ;
        RECT  2.690 1.370 3.480 1.610 ;
        RECT  2.690 1.020 2.930 1.610 ;
        RECT  2.370 3.940 2.870 4.340 ;
        RECT  2.630 2.930 2.870 4.340 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  5.600 3.060 6.000 5.600 ;
        RECT  4.230 2.780 4.630 5.600 ;
        RECT  3.110 4.180 3.510 5.600 ;
        RECT  1.320 4.620 1.720 5.600 ;
        RECT  0.150 3.050 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.830 0.000 5.230 0.980 ;
        RECT  3.350 0.000 3.750 0.980 ;
        RECT  1.850 0.000 2.250 0.980 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.100 1.370 1.340 ;
        RECT  1.130 1.100 1.370 1.710 ;
        RECT  1.130 1.470 2.170 1.710 ;
        RECT  1.930 1.850 2.990 2.250 ;
        RECT  1.930 1.470 2.170 3.440 ;
        RECT  0.800 3.200 2.170 3.440 ;
        RECT  0.800 3.200 1.040 4.140 ;
    END
END an02d7

MACRO an02d4
    CLASS CORE ;
    FOREIGN an02d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.397  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.470 0.500 3.020 ;
        RECT  0.220 1.890 0.460 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.980 2.520 1.620 3.020 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.179  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.060 3.740 3.690 4.140 ;
        RECT  3.450 1.450 3.690 4.140 ;
        RECT  1.960 1.450 3.690 1.690 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.920 5.600 ;
        RECT  2.800 4.610 3.200 5.600 ;
        RECT  1.500 4.610 1.900 5.600 ;
        RECT  0.230 4.030 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.920 0.740 ;
        RECT  2.750 0.000 3.150 0.970 ;
        RECT  1.370 0.000 1.780 0.930 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.170 1.720 1.410 ;
        RECT  1.480 1.170 1.720 2.230 ;
        RECT  1.480 1.990 2.100 2.230 ;
        RECT  1.860 2.320 2.970 2.720 ;
        RECT  1.860 1.990 2.100 3.500 ;
        RECT  0.730 3.260 2.100 3.500 ;
    END
END an02d4

MACRO an02d2
    CLASS CORE ;
    FOREIGN an02d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.252  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.460 0.500 3.020 ;
        RECT  0.220 1.890 0.460 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.252  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.980 2.520 1.620 3.020 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.663  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.740 2.580 4.140 ;
        RECT  2.340 1.450 2.580 4.140 ;
        RECT  1.960 1.450 2.580 1.690 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 3.360 5.600 ;
        RECT  2.890 4.140 3.130 5.600 ;
        RECT  1.390 4.360 1.630 5.600 ;
        RECT  0.230 4.070 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 3.360 0.740 ;
        RECT  2.890 0.000 3.130 1.150 ;
        RECT  1.370 0.000 1.780 0.930 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.170 1.720 1.410 ;
        RECT  1.480 1.170 1.720 2.280 ;
        RECT  1.480 2.040 2.100 2.280 ;
        RECT  1.860 2.040 2.100 3.500 ;
        RECT  0.740 3.260 2.100 3.500 ;
    END
END an02d2

MACRO an02d1
    CLASS CORE ;
    FOREIGN an02d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.080 0.800 2.450 ;
        RECT  0.120 2.080 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.080 2.020 1.620 2.520 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.473  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.200 2.680 4.140 ;
        RECT  2.340 1.050 2.680 4.140 ;
        RECT  2.330 1.050 2.680 1.450 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  1.440 4.250 1.680 5.600 ;
        RECT  0.230 4.250 0.470 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  1.400 0.000 1.800 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 2.100 1.780 ;
        RECT  1.860 1.540 2.100 3.010 ;
        RECT  0.820 2.770 2.100 3.010 ;
        RECT  0.820 2.770 1.060 3.450 ;
    END
END an02d1

MACRO an02d0
    CLASS CORE ;
    FOREIGN an02d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.080 0.800 2.450 ;
        RECT  0.120 2.080 0.500 3.020 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.080 2.020 1.620 2.520 ;
        END
    END A2
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.913  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 3.200 2.680 4.140 ;
        RECT  2.340 1.050 2.680 4.140 ;
        RECT  2.330 1.050 2.680 1.450 ;
        END
    END Z
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 2.800 5.600 ;
        RECT  1.140 4.700 1.560 5.600 ;
        RECT  0.150 4.710 0.550 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 2.800 0.740 ;
        RECT  1.400 0.000 1.800 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.540 2.100 1.780 ;
        RECT  1.860 1.540 2.100 3.010 ;
        RECT  0.820 2.770 2.100 3.010 ;
        RECT  0.820 2.770 1.060 3.450 ;
    END
END an02d0

MACRO ah01d4
    CLASS CORE ;
    FOREIGN ah01d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.402  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.830 1.430 6.660 1.990 ;
        RECT  5.830 1.380 6.220 1.990 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.748  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.500 2.520 4.980 3.070 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.802  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.410 2.020 8.840 2.460 ;
        RECT  8.420 1.070 8.810 1.500 ;
        RECT  6.800 3.400 8.650 3.640 ;
        RECT  8.410 1.220 8.650 3.640 ;
        RECT  6.920 1.220 8.810 1.460 ;
        RECT  6.920 1.070 7.320 1.470 ;
        RECT  6.800 3.400 7.040 4.620 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.230 3.050 2.600 3.470 ;
        RECT  0.230 1.770 1.120 2.170 ;
        RECT  0.230 1.770 0.500 3.470 ;
        RECT  0.120 2.580 0.500 3.020 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 8.960 5.600 ;
        RECT  7.720 3.880 7.960 5.600 ;
        RECT  6.060 3.030 6.300 5.600 ;
        RECT  4.490 4.560 4.930 5.600 ;
        RECT  2.840 4.060 3.080 5.600 ;
        RECT  1.540 3.810 1.780 5.600 ;
        RECT  0.240 3.820 0.480 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 8.960 0.740 ;
        RECT  7.690 0.000 8.090 0.980 ;
        RECT  6.180 0.000 6.580 0.980 ;
        RECT  3.390 0.000 3.790 0.980 ;
        RECT  1.540 0.000 1.780 1.930 ;
        RECT  0.230 0.000 0.470 1.450 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  4.550 1.480 5.110 1.720 ;
        RECT  4.550 1.480 4.790 2.240 ;
        RECT  4.020 2.000 4.790 2.240 ;
        RECT  0.740 2.410 3.080 2.810 ;
        RECT  2.840 2.410 3.080 3.530 ;
        RECT  4.020 2.000 4.260 3.530 ;
        RECT  2.840 3.290 4.260 3.530 ;
        RECT  4.070 0.980 5.590 1.220 ;
        RECT  4.070 0.980 4.310 1.760 ;
        RECT  2.160 1.520 4.310 1.760 ;
        RECT  5.350 0.980 5.590 2.560 ;
        RECT  5.120 1.960 5.590 2.320 ;
        RECT  7.670 1.840 7.910 2.560 ;
        RECT  5.220 2.320 7.910 2.560 ;
        RECT  3.320 1.520 3.560 2.920 ;
        RECT  5.220 1.960 5.460 3.540 ;
        RECT  5.420 3.300 5.660 4.040 ;
    END
END ah01d4

MACRO ah01d2
    CLASS CORE ;
    FOREIGN ah01d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 2.370 3.740 3.770 ;
        RECT  0.630 2.370 3.740 2.610 ;
        RECT  0.630 1.730 1.060 2.610 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.700 1.460 2.100 2.130 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.164  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.220 2.580 6.850 3.020 ;
        RECT  6.610 1.550 6.850 3.020 ;
        RECT  6.440 2.580 6.680 3.870 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.172  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.130 1.550 5.380 3.870 ;
        RECT  4.530 2.100 5.380 2.380 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 7.840 5.600 ;
        RECT  7.180 4.480 7.420 5.600 ;
        RECT  5.880 4.480 6.120 5.600 ;
        RECT  4.570 4.480 4.810 5.600 ;
        RECT  2.470 4.620 2.870 5.600 ;
        RECT  0.980 4.040 1.220 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 7.840 0.740 ;
        RECT  7.350 0.000 7.590 1.420 ;
        RECT  5.870 0.000 6.110 1.420 ;
        RECT  4.390 0.000 4.630 1.420 ;
        RECT  3.540 0.000 3.940 0.980 ;
        RECT  1.750 0.000 1.990 1.200 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.060 0.550 1.380 ;
        RECT  0.150 1.060 0.390 3.610 ;
        RECT  0.150 3.290 2.600 3.610 ;
        RECT  3.100 1.730 4.220 2.050 ;
        RECT  3.980 2.950 4.500 3.350 ;
        RECT  1.700 4.140 4.220 4.380 ;
        RECT  3.980 1.730 4.220 4.460 ;
        RECT  3.700 4.140 4.220 4.460 ;
    END
END ah01d2

MACRO ah01d1
    CLASS CORE ;
    FOREIGN ah01d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.200 2.810 3.440 3.380 ;
        RECT  0.630 2.810 3.440 3.050 ;
        RECT  0.630 2.440 0.980 3.050 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.750 2.180 2.460 ;
        RECT  1.080 1.750 2.180 2.150 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.053  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.610 2.580 6.040 3.870 ;
        RECT  5.800 1.550 6.040 3.870 ;
        RECT  5.460 1.550 6.040 1.950 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.036  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.400 2.020 4.980 2.460 ;
        RECT  4.310 3.550 4.690 3.870 ;
        RECT  4.400 1.620 4.690 3.870 ;
        RECT  4.010 1.620 4.690 1.860 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.160 5.600 ;
        RECT  4.960 4.480 5.200 5.600 ;
        RECT  2.410 4.620 2.810 5.600 ;
        RECT  0.920 4.140 1.160 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.160 0.740 ;
        RECT  4.830 0.000 5.070 1.420 ;
        RECT  3.130 0.000 3.530 0.980 ;
        RECT  1.430 0.000 1.670 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.220 0.550 1.540 ;
        RECT  0.150 1.220 0.390 3.610 ;
        RECT  0.150 3.290 2.600 3.610 ;
        RECT  2.690 1.750 3.760 2.150 ;
        RECT  3.520 1.750 3.760 2.430 ;
        RECT  3.720 2.950 4.160 3.350 ;
        RECT  3.720 2.190 3.960 4.460 ;
        RECT  1.640 4.140 4.010 4.380 ;
        RECT  3.720 4.050 4.010 4.460 ;
        RECT  3.590 4.140 4.010 4.460 ;
    END
END ah01d1

MACRO ah01d0
    CLASS CORE ;
    FOREIGN ah01d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.490 2.390 3.730 3.770 ;
        RECT  0.630 2.390 3.730 2.630 ;
        RECT  0.630 2.020 1.060 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.340 1.460 2.180 1.900 ;
        RECT  1.340 1.460 1.740 2.150 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.598  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.930 1.460 6.170 3.710 ;
        RECT  5.660 2.580 6.170 3.020 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.598  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.450 2.580 4.980 3.020 ;
        RECT  4.450 1.750 4.690 3.710 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 6.720 5.600 ;
        RECT  5.190 3.610 5.430 5.600 ;
        RECT  2.310 4.620 2.710 5.600 ;
        RECT  0.820 3.940 1.060 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 6.720 0.740 ;
        RECT  5.190 0.000 5.430 2.090 ;
        RECT  3.540 0.000 3.940 0.980 ;
        RECT  1.750 0.000 1.990 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.150 1.220 0.550 1.540 ;
        RECT  0.150 1.220 0.390 3.450 ;
        RECT  2.350 2.950 2.750 3.450 ;
        RECT  0.150 3.130 2.750 3.450 ;
        RECT  3.810 1.410 4.050 2.090 ;
        RECT  3.100 1.850 4.210 2.090 ;
        RECT  3.970 1.850 4.210 4.460 ;
        RECT  1.540 4.140 4.210 4.380 ;
        RECT  3.660 4.220 4.950 4.460 ;
        RECT  1.540 4.140 1.860 4.560 ;
    END
END ah01d0

MACRO adp1d4
    CLASS CORE ;
    FOREIGN adp1d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.379  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 2.580 0.540 3.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.051  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.820 2.450 5.030 2.690 ;
        RECT  3.820 1.130 4.060 2.690 ;
        RECT  2.860 1.130 4.060 1.370 ;
        RECT  2.180 1.520 3.100 1.760 ;
        RECT  2.860 1.130 3.100 1.760 ;
        RECT  2.180 1.520 2.420 2.640 ;
        RECT  1.740 2.400 2.180 3.020 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.666  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.580 2.660 10.360 2.900 ;
        RECT  9.580 2.480 10.040 3.020 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.921  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.190 1.360 20.010 1.600 ;
        RECT  19.300 1.360 19.540 4.380 ;
        RECT  18.810 4.380 19.370 4.620 ;
        RECT  19.130 4.140 19.540 4.380 ;
        RECT  17.690 2.980 19.540 3.220 ;
        RECT  19.100 1.360 19.540 3.220 ;
        END
    END CO
    PIN P
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.209  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.090 1.010 14.650 1.250 ;
        RECT  13.090 1.220 14.330 1.460 ;
        RECT  12.940 2.370 14.060 3.050 ;
        RECT  13.700 1.220 14.060 3.050 ;
        RECT  12.770 1.000 13.330 1.240 ;
        RECT  12.100 2.760 14.060 3.000 ;
        END
    END P
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.941  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.520 1.360 17.220 1.600 ;
        RECT  14.940 3.130 16.790 3.580 ;
        RECT  16.370 1.360 16.790 3.580 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 20.160 5.600 ;
        RECT  19.610 4.620 20.010 5.600 ;
        RECT  17.770 3.600 18.650 4.000 ;
        RECT  17.770 3.600 18.170 5.600 ;
        RECT  16.950 4.620 17.350 5.600 ;
        RECT  15.650 4.620 16.050 5.600 ;
        RECT  14.160 4.620 14.560 5.600 ;
        RECT  12.860 4.620 13.260 5.600 ;
        RECT  10.770 4.710 11.170 5.600 ;
        RECT  9.470 4.710 9.870 5.600 ;
        RECT  7.170 4.710 7.570 5.600 ;
        RECT  4.290 4.710 4.690 5.600 ;
        RECT  1.990 4.380 2.390 5.600 ;
        RECT  0.720 4.320 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 20.160 0.740 ;
        RECT  19.000 0.000 19.400 0.980 ;
        RECT  17.630 0.000 18.030 0.980 ;
        RECT  16.260 0.000 16.660 0.980 ;
        RECT  15.000 0.000 15.390 0.980 ;
        RECT  13.570 0.000 13.850 0.980 ;
        RECT  12.000 0.000 12.400 0.890 ;
        RECT  10.030 0.000 10.430 0.890 ;
        RECT  9.230 0.000 9.630 1.260 ;
        RECT  6.770 0.000 7.170 1.260 ;
        RECT  4.490 0.000 4.890 0.890 ;
        RECT  2.320 0.000 2.620 1.280 ;
        RECT  0.630 0.000 1.030 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.260 0.980 2.080 1.220 ;
        RECT  1.260 1.850 1.910 2.090 ;
        RECT  1.260 0.980 1.500 3.600 ;
        RECT  1.260 3.360 1.860 3.600 ;
        RECT  0.150 1.850 1.020 2.090 ;
        RECT  0.780 1.850 1.020 4.080 ;
        RECT  0.150 3.720 1.020 3.960 ;
        RECT  0.760 3.840 1.700 4.080 ;
        RECT  1.530 3.900 2.870 4.140 ;
        RECT  2.630 3.900 2.870 4.620 ;
        RECT  2.630 4.380 3.950 4.620 ;
        RECT  5.100 4.380 6.800 4.620 ;
        RECT  9.040 1.980 10.130 2.220 ;
        RECT  6.940 2.460 7.500 2.700 ;
        RECT  7.260 2.460 7.500 3.180 ;
        RECT  9.040 1.980 9.280 3.180 ;
        RECT  7.260 2.940 9.340 3.180 ;
        RECT  9.090 2.940 9.340 3.510 ;
        RECT  9.090 3.270 10.370 3.510 ;
        RECT  11.120 1.770 11.500 2.000 ;
        RECT  11.120 1.520 11.440 2.000 ;
        RECT  11.260 1.840 11.770 2.060 ;
        RECT  11.330 1.840 11.770 2.450 ;
        RECT  11.330 1.840 11.570 3.010 ;
        RECT  11.140 2.770 11.380 3.500 ;
        RECT  11.140 3.260 11.700 3.500 ;
        RECT  5.060 1.060 6.470 1.220 ;
        RECT  11.680 1.110 11.860 1.590 ;
        RECT  5.120 0.980 6.470 1.220 ;
        RECT  7.410 0.980 8.800 1.220 ;
        RECT  10.660 1.040 11.800 1.280 ;
        RECT  4.580 1.130 5.350 1.330 ;
        RECT  11.620 1.160 11.920 1.340 ;
        RECT  11.680 1.160 11.920 1.590 ;
        RECT  4.580 1.130 5.310 1.370 ;
        RECT  10.530 1.130 10.890 1.370 ;
        RECT  6.230 0.980 6.470 1.740 ;
        RECT  11.680 1.350 12.420 1.590 ;
        RECT  12.160 1.350 12.420 2.080 ;
        RECT  7.410 0.980 7.650 1.740 ;
        RECT  6.230 1.500 7.650 1.740 ;
        RECT  8.560 1.500 10.770 1.740 ;
        RECT  4.580 1.130 4.820 2.210 ;
        RECT  4.580 2.000 5.400 2.210 ;
        RECT  12.160 1.700 13.460 2.080 ;
        RECT  4.580 1.970 5.350 2.210 ;
        RECT  10.530 1.130 10.770 2.480 ;
        RECT  5.200 2.040 5.510 2.270 ;
        RECT  3.340 1.610 3.580 2.430 ;
        RECT  10.530 2.240 11.090 2.480 ;
        RECT  8.560 0.980 8.800 2.700 ;
        RECT  7.830 2.460 8.800 2.700 ;
        RECT  5.270 2.040 5.510 3.170 ;
        RECT  3.270 2.930 5.510 3.170 ;
        RECT  3.270 2.250 3.510 4.020 ;
        RECT  8.080 1.460 8.320 2.220 ;
        RECT  6.460 1.980 8.320 2.220 ;
        RECT  14.300 1.890 15.760 2.290 ;
        RECT  6.460 1.980 6.700 3.660 ;
        RECT  14.300 1.890 14.540 3.530 ;
        RECT  11.940 3.290 14.540 3.530 ;
        RECT  6.460 3.420 8.800 3.660 ;
        RECT  8.560 3.420 8.800 3.990 ;
        RECT  11.940 3.290 12.180 3.990 ;
        RECT  8.560 3.750 12.180 3.990 ;
        RECT  5.540 1.480 5.990 1.800 ;
        RECT  5.620 1.480 5.990 1.820 ;
        RECT  17.050 2.330 18.380 2.730 ;
        RECT  5.750 1.480 5.990 4.140 ;
        RECT  5.740 3.280 5.990 4.140 ;
        RECT  5.740 3.900 7.330 4.140 ;
        RECT  7.090 3.900 7.330 4.470 ;
        RECT  12.450 4.140 17.290 4.380 ;
        RECT  17.050 2.330 17.290 4.380 ;
        RECT  7.090 4.230 12.660 4.470 ;
    END
END adp1d4

MACRO adp1d2
    CLASS CORE ;
    FOREIGN adp1d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.292  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.700 2.640 11.470 3.020 ;
        RECT  11.070 2.360 11.470 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.020 2.570 9.930 2.940 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.733  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.830 1.880 12.070 2.670 ;
        RECT  11.060 1.880 12.070 2.120 ;
        RECT  11.060 1.140 11.300 2.120 ;
        RECT  8.200 1.140 11.300 1.380 ;
        RECT  1.220 1.220 8.420 1.460 ;
        RECT  0.140 1.130 1.480 1.370 ;
        RECT  0.140 2.440 0.500 3.360 ;
        RECT  0.140 1.130 0.380 3.360 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.086  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.530 3.460 15.000 3.780 ;
        RECT  14.760 1.700 15.000 3.780 ;
        RECT  14.530 1.700 15.000 2.460 ;
        END
    END CO
    PIN P
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.378  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.710 1.700 6.110 2.380 ;
        RECT  5.380 2.220 5.750 2.490 ;
        RECT  5.570 2.100 6.110 2.380 ;
        RECT  5.380 2.220 5.620 3.580 ;
        END
    END P
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.989  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 3.140 1.840 3.580 ;
        RECT  1.220 1.700 1.680 2.030 ;
        RECT  1.220 1.700 1.460 3.580 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.680 5.600 ;
        RECT  14.050 4.150 14.290 5.600 ;
        RECT  11.000 4.620 11.400 5.600 ;
        RECT  9.800 4.620 10.200 5.600 ;
        RECT  8.680 4.620 9.080 5.600 ;
        RECT  6.410 4.300 6.650 5.600 ;
        RECT  4.370 4.300 4.610 5.600 ;
        RECT  2.040 4.300 2.280 5.600 ;
        RECT  0.500 4.300 0.740 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.680 0.740 ;
        RECT  13.950 0.000 14.350 0.980 ;
        RECT  11.540 0.000 11.780 1.640 ;
        RECT  9.010 0.000 9.410 0.890 ;
        RECT  6.390 0.000 6.790 0.980 ;
        RECT  5.000 0.000 5.400 0.970 ;
        RECT  4.160 0.000 4.560 0.980 ;
        RECT  1.880 0.000 2.280 0.890 ;
        RECT  0.510 0.000 0.910 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.500 1.760 3.510 2.000 ;
        RECT  1.700 2.650 2.740 2.890 ;
        RECT  2.500 1.760 2.740 3.580 ;
        RECT  2.500 3.340 3.560 3.580 ;
        RECT  0.620 1.610 0.860 2.230 ;
        RECT  0.740 2.020 0.980 4.060 ;
        RECT  0.640 3.560 0.980 4.060 ;
        RECT  4.170 2.730 4.410 4.060 ;
        RECT  0.640 3.820 4.410 4.060 ;
        RECT  6.750 1.700 8.020 1.940 ;
        RECT  5.960 2.620 6.990 2.860 ;
        RECT  6.750 1.700 6.990 3.510 ;
        RECT  6.750 3.270 7.800 3.510 ;
        RECT  8.520 1.680 10.200 1.920 ;
        RECT  8.110 2.300 8.760 2.540 ;
        RECT  8.520 1.680 8.760 3.420 ;
        RECT  8.520 3.180 9.680 3.420 ;
        RECT  10.580 1.700 10.820 2.400 ;
        RECT  10.220 2.160 10.820 2.400 ;
        RECT  7.450 2.280 7.690 3.030 ;
        RECT  7.450 2.790 8.280 3.030 ;
        RECT  10.220 3.280 11.040 3.520 ;
        RECT  8.040 2.790 8.280 3.900 ;
        RECT  10.220 2.160 10.460 3.900 ;
        RECT  8.040 3.660 10.460 3.900 ;
        RECT  4.770 1.700 5.330 1.940 ;
        RECT  4.770 1.700 5.010 2.480 ;
        RECT  2.990 2.240 5.140 2.480 ;
        RECT  2.990 2.240 3.230 3.000 ;
        RECT  12.000 2.910 13.100 3.150 ;
        RECT  12.000 2.910 12.240 3.500 ;
        RECT  11.280 3.260 12.240 3.500 ;
        RECT  4.900 2.240 5.140 4.570 ;
        RECT  4.900 3.820 7.130 4.060 ;
        RECT  6.890 3.820 7.130 4.380 ;
        RECT  11.280 3.260 11.520 4.380 ;
        RECT  6.890 4.140 11.520 4.380 ;
        RECT  4.900 3.820 5.460 4.570 ;
        RECT  11.930 4.190 13.630 4.430 ;
        RECT  12.680 1.320 14.290 1.560 ;
        RECT  14.050 2.830 14.460 3.230 ;
        RECT  14.050 1.320 14.290 3.680 ;
        RECT  12.490 3.440 14.290 3.680 ;
    END
END adp1d2

MACRO adp1d1
    CLASS CORE ;
    FOREIGN adp1d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.286  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.120 2.360 11.620 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.470 2.570 10.020 2.940 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.727  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.880 1.880 12.120 2.670 ;
        RECT  11.110 1.880 12.120 2.120 ;
        RECT  11.110 1.220 11.350 2.120 ;
        RECT  1.220 1.220 11.350 1.460 ;
        RECT  0.140 1.130 1.480 1.370 ;
        RECT  0.140 2.440 0.540 3.340 ;
        RECT  0.140 1.130 0.380 3.340 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.143  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.570 3.460 15.000 3.780 ;
        RECT  14.760 1.700 15.000 3.780 ;
        RECT  14.550 1.700 15.000 2.460 ;
        END
    END CO
    PIN P
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.378  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.760 1.700 6.100 2.380 ;
        RECT  5.570 2.100 6.100 2.380 ;
        RECT  5.380 2.220 5.750 2.490 ;
        RECT  5.380 2.220 5.620 3.580 ;
        END
    END P
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.989  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 3.140 1.790 3.580 ;
        RECT  1.260 1.700 1.730 2.030 ;
        RECT  1.260 1.700 1.500 3.580 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.120 5.600 ;
        RECT  14.050 4.190 14.290 5.600 ;
        RECT  11.140 4.620 11.560 5.600 ;
        RECT  9.800 4.620 10.200 5.600 ;
        RECT  8.680 4.620 9.080 5.600 ;
        RECT  6.410 4.300 6.650 5.600 ;
        RECT  4.370 4.300 4.610 5.600 ;
        RECT  2.040 4.300 2.280 5.600 ;
        RECT  0.500 4.300 0.740 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.120 0.740 ;
        RECT  14.000 0.000 14.410 0.980 ;
        RECT  11.590 0.000 11.830 1.640 ;
        RECT  9.060 0.000 9.460 0.890 ;
        RECT  6.440 0.000 6.840 0.980 ;
        RECT  4.210 0.000 4.610 0.980 ;
        RECT  1.930 0.000 2.330 0.890 ;
        RECT  0.560 0.000 0.960 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.500 1.760 3.560 2.000 ;
        RECT  1.740 2.360 2.740 2.600 ;
        RECT  2.500 1.760 2.740 3.580 ;
        RECT  2.500 3.340 3.560 3.580 ;
        RECT  0.670 1.610 0.910 2.230 ;
        RECT  0.780 2.020 1.020 4.060 ;
        RECT  0.640 3.560 1.020 4.060 ;
        RECT  4.170 2.730 4.410 4.060 ;
        RECT  0.640 3.820 4.410 4.060 ;
        RECT  6.920 1.700 8.070 1.940 ;
        RECT  5.960 2.620 7.160 2.860 ;
        RECT  6.920 1.700 7.160 3.510 ;
        RECT  6.920 3.270 7.850 3.510 ;
        RECT  8.570 1.700 10.250 1.940 ;
        RECT  8.160 2.230 8.810 2.470 ;
        RECT  8.570 1.700 8.810 3.420 ;
        RECT  8.570 3.180 9.680 3.420 ;
        RECT  10.630 1.700 10.870 2.450 ;
        RECT  10.330 2.210 10.870 2.450 ;
        RECT  7.500 2.280 7.740 3.030 ;
        RECT  7.500 2.790 8.330 3.030 ;
        RECT  10.330 3.280 11.040 3.520 ;
        RECT  8.090 2.790 8.330 3.900 ;
        RECT  10.330 2.210 10.570 3.900 ;
        RECT  8.090 3.660 10.570 3.900 ;
        RECT  4.830 1.700 5.380 1.940 ;
        RECT  4.830 1.700 5.070 2.480 ;
        RECT  2.990 2.240 5.140 2.480 ;
        RECT  2.990 2.240 3.230 3.000 ;
        RECT  12.000 2.910 13.100 3.150 ;
        RECT  12.000 2.910 12.240 3.500 ;
        RECT  11.280 3.260 12.240 3.500 ;
        RECT  4.900 2.240 5.140 4.570 ;
        RECT  4.900 3.820 7.130 4.060 ;
        RECT  6.890 3.820 7.130 4.380 ;
        RECT  11.280 3.260 11.520 4.380 ;
        RECT  6.890 4.140 11.520 4.380 ;
        RECT  4.900 3.820 5.460 4.570 ;
        RECT  11.930 4.190 13.630 4.430 ;
        RECT  12.730 1.320 14.310 1.560 ;
        RECT  14.070 2.830 14.490 3.230 ;
        RECT  14.070 1.320 14.310 3.680 ;
        RECT  12.490 3.440 14.310 3.680 ;
    END
END adp1d1

MACRO adp1d0
    CLASS CORE ;
    FOREIGN adp1d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.120 2.360 11.620 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.470 2.570 10.020 2.940 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.736  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.880 1.880 12.120 2.670 ;
        RECT  11.110 1.880 12.120 2.120 ;
        RECT  11.110 1.220 11.350 2.120 ;
        RECT  1.220 1.220 11.350 1.460 ;
        RECT  0.140 1.130 1.480 1.370 ;
        RECT  0.140 2.580 0.540 3.330 ;
        RECT  0.140 1.130 0.380 3.330 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.697  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.560 3.440 15.000 3.760 ;
        RECT  14.760 1.700 15.000 3.760 ;
        RECT  14.550 1.700 15.000 2.460 ;
        END
    END CO
    PIN P
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.374  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.760 1.700 6.100 2.380 ;
        RECT  5.570 2.100 6.100 2.380 ;
        RECT  5.360 2.220 5.750 2.470 ;
        RECT  5.360 2.220 5.600 3.580 ;
        END
    END P
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.989  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 3.140 1.770 3.580 ;
        RECT  1.260 1.700 1.730 2.030 ;
        RECT  1.260 1.700 1.500 3.580 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.120 5.600 ;
        RECT  14.040 4.180 14.280 5.600 ;
        RECT  11.100 4.620 11.520 5.600 ;
        RECT  9.790 4.620 10.190 5.600 ;
        RECT  8.660 4.620 9.060 5.600 ;
        RECT  6.390 4.300 6.630 5.600 ;
        RECT  4.350 4.300 4.590 5.600 ;
        RECT  2.020 4.300 2.260 5.600 ;
        RECT  0.500 4.300 0.740 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.120 0.740 ;
        RECT  14.000 0.000 14.400 0.980 ;
        RECT  11.590 0.000 11.830 1.640 ;
        RECT  9.060 0.000 9.460 0.890 ;
        RECT  6.440 0.000 6.840 0.980 ;
        RECT  5.040 0.000 5.440 0.970 ;
        RECT  4.210 0.000 4.610 0.980 ;
        RECT  1.930 0.000 2.330 0.890 ;
        RECT  0.560 0.000 0.960 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.500 1.760 3.560 2.000 ;
        RECT  1.740 2.360 2.740 2.600 ;
        RECT  2.500 1.760 2.740 3.580 ;
        RECT  2.500 3.340 3.540 3.580 ;
        RECT  0.670 1.610 0.910 2.320 ;
        RECT  0.780 2.030 1.020 4.060 ;
        RECT  0.620 3.560 1.020 4.060 ;
        RECT  4.170 2.730 4.410 4.060 ;
        RECT  0.620 3.820 4.410 4.060 ;
        RECT  6.920 1.700 8.070 1.940 ;
        RECT  5.940 2.620 7.160 2.860 ;
        RECT  6.920 1.700 7.160 3.510 ;
        RECT  6.920 3.270 7.830 3.510 ;
        RECT  8.570 1.700 10.250 1.940 ;
        RECT  8.140 2.230 8.810 2.470 ;
        RECT  8.570 1.700 8.810 3.420 ;
        RECT  8.570 3.180 9.660 3.420 ;
        RECT  10.630 1.700 10.870 2.450 ;
        RECT  10.330 2.210 10.870 2.450 ;
        RECT  7.500 2.280 7.740 3.030 ;
        RECT  7.500 2.790 8.330 3.030 ;
        RECT  10.330 3.280 11.040 3.520 ;
        RECT  8.090 2.790 8.330 3.900 ;
        RECT  10.330 2.210 10.570 3.900 ;
        RECT  8.090 3.660 10.570 3.900 ;
        RECT  4.830 1.700 5.380 1.940 ;
        RECT  4.830 1.700 5.070 2.480 ;
        RECT  2.990 2.240 5.120 2.480 ;
        RECT  2.990 2.240 3.230 3.000 ;
        RECT  11.970 2.910 13.100 3.150 ;
        RECT  11.970 2.910 12.210 3.500 ;
        RECT  11.280 3.260 12.210 3.500 ;
        RECT  4.880 2.240 5.120 4.570 ;
        RECT  4.880 3.820 7.130 4.060 ;
        RECT  6.890 3.820 7.130 4.380 ;
        RECT  11.280 3.260 11.520 4.380 ;
        RECT  6.890 4.140 11.520 4.380 ;
        RECT  4.880 3.820 5.460 4.570 ;
        RECT  11.890 4.260 13.590 4.500 ;
        RECT  12.730 1.320 14.310 1.560 ;
        RECT  14.070 2.810 14.480 3.210 ;
        RECT  14.070 1.320 14.310 3.680 ;
        RECT  12.450 3.440 14.310 3.680 ;
    END
END adp1d0

MACRO adiode
    CLASS CORE ;
    FOREIGN adiode 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNADIFFAREA 0.925  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.560 3.450 ;
        END
    END I
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 1.120 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 1.120 0.740 ;
        END
    END VSS
END adiode

MACRO ad01d4
    CLASS CORE ;
    FOREIGN ad01d4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.451  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.380 2.020 2.360 2.460 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.583  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.320 1.670 6.560 2.600 ;
        RECT  5.690 1.670 6.560 1.910 ;
        RECT  5.690 0.990 5.930 1.910 ;
        RECT  3.480 0.990 5.930 1.230 ;
        RECT  2.600 2.020 3.720 2.460 ;
        RECT  3.480 0.990 3.720 2.460 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.420  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.560 1.060 3.040 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.963  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.490 1.970 11.730 4.150 ;
        RECT  10.000 1.730 11.720 1.970 ;
        RECT  10.180 3.220 11.730 3.460 ;
        RECT  11.480 0.980 11.720 3.460 ;
        RECT  11.260 1.970 11.730 3.460 ;
        RECT  10.180 3.220 10.420 3.920 ;
        RECT  10.000 1.110 10.240 1.970 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.051  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.960 1.430 14.680 1.670 ;
        RECT  14.440 0.980 14.680 1.670 ;
        RECT  12.790 2.580 14.500 2.970 ;
        RECT  14.060 1.430 14.500 2.970 ;
        RECT  12.960 0.980 13.200 1.670 ;
        RECT  12.790 2.580 13.030 4.340 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 15.120 5.600 ;
        RECT  14.620 4.310 14.860 5.600 ;
        RECT  13.350 3.260 13.590 5.600 ;
        RECT  12.150 4.620 12.550 5.600 ;
        RECT  10.850 4.620 11.250 5.600 ;
        RECT  9.530 4.620 9.930 5.600 ;
        RECT  7.540 4.700 7.940 5.600 ;
        RECT  6.150 4.700 6.550 5.600 ;
        RECT  2.810 4.400 3.050 5.600 ;
        RECT  1.500 4.400 1.740 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 15.120 0.740 ;
        RECT  13.700 0.000 13.940 1.150 ;
        RECT  12.220 0.000 12.460 1.380 ;
        RECT  10.740 0.000 10.980 1.200 ;
        RECT  7.690 0.000 8.090 0.890 ;
        RECT  6.510 0.000 6.910 0.890 ;
        RECT  3.000 0.000 3.240 1.770 ;
        RECT  1.340 0.000 1.740 0.910 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 3.330 2.400 3.570 ;
        RECT  0.870 1.300 2.580 1.540 ;
        RECT  7.390 3.000 8.640 3.240 ;
        RECT  7.390 3.000 7.630 3.610 ;
        RECT  6.870 3.370 7.630 3.610 ;
        RECT  7.100 1.630 8.860 1.870 ;
        RECT  9.470 0.980 9.710 1.730 ;
        RECT  9.280 1.490 9.520 2.320 ;
        RECT  6.910 2.110 9.400 2.350 ;
        RECT  6.910 2.110 7.150 3.080 ;
        RECT  4.900 2.840 7.150 3.080 ;
        RECT  9.160 2.110 9.400 3.890 ;
        RECT  8.830 3.650 9.400 3.890 ;
        RECT  4.900 1.470 5.140 4.110 ;
        RECT  4.490 3.870 5.140 4.110 ;
        RECT  3.960 1.520 4.520 1.760 ;
        RECT  0.230 1.210 0.470 2.000 ;
        RECT  9.800 2.270 10.750 2.690 ;
        RECT  3.120 3.240 4.200 3.560 ;
        RECT  3.960 1.520 4.200 3.640 ;
        RECT  3.790 3.240 4.200 3.640 ;
        RECT  0.120 1.770 0.360 4.050 ;
        RECT  3.120 3.240 3.370 4.050 ;
        RECT  0.120 3.810 3.370 4.050 ;
        RECT  3.870 3.240 4.110 4.620 ;
        RECT  5.380 4.140 9.940 4.380 ;
        RECT  9.700 2.480 9.940 4.380 ;
        RECT  0.230 3.810 0.470 4.610 ;
        RECT  3.870 4.380 5.620 4.620 ;
    END
END ad01d4

MACRO ad01d2
    CLASS CORE ;
    FOREIGN ad01d2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.802  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.630 7.440 2.870 ;
        RECT  7.200 2.100 7.440 2.870 ;
        RECT  2.860 2.630 3.300 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.637  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.120 2.020 3.860 2.390 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.020  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.980 2.100 6.840 2.390 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.181  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.160 1.770 10.580 3.650 ;
        RECT  10.050 1.770 10.580 2.100 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.284  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.580 3.330 9.220 3.570 ;
        RECT  8.970 2.220 9.220 3.570 ;
        RECT  8.460 2.020 9.010 2.460 ;
        RECT  8.770 1.570 9.010 2.460 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 11.200 5.600 ;
        RECT  10.730 4.280 10.970 5.600 ;
        RECT  9.420 4.290 9.660 5.600 ;
        RECT  8.090 4.290 8.330 5.600 ;
        RECT  4.700 4.700 5.120 5.600 ;
        RECT  3.450 4.140 3.690 5.600 ;
        RECT  0.850 4.140 1.090 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 11.200 0.740 ;
        RECT  10.650 0.000 11.050 0.890 ;
        RECT  9.460 0.000 9.860 0.890 ;
        RECT  7.950 0.000 8.190 1.280 ;
        RECT  4.870 0.000 5.110 1.280 ;
        RECT  3.450 0.000 3.690 1.340 ;
        RECT  0.820 0.000 1.060 1.270 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.170 1.630 1.880 1.870 ;
        RECT  0.150 3.600 1.910 3.840 ;
        RECT  4.040 1.620 5.820 1.860 ;
        RECT  4.360 3.130 6.060 3.370 ;
        RECT  5.820 3.130 6.060 4.120 ;
        RECT  6.180 0.980 6.420 1.840 ;
        RECT  6.180 1.600 8.110 1.840 ;
        RECT  7.870 2.800 8.700 3.040 ;
        RECT  7.870 1.600 8.110 3.370 ;
        RECT  6.310 3.130 8.110 3.370 ;
        RECT  2.250 0.980 2.490 2.350 ;
        RECT  0.120 2.110 2.490 2.350 ;
        RECT  0.120 2.110 0.360 3.360 ;
        RECT  0.120 3.120 2.480 3.360 ;
        RECT  2.240 3.660 5.580 3.900 ;
        RECT  9.680 2.390 9.920 4.050 ;
        RECT  6.390 3.810 9.920 4.050 ;
        RECT  5.340 3.660 5.580 4.600 ;
        RECT  2.240 3.120 2.480 4.540 ;
        RECT  5.340 4.360 6.630 4.600 ;
        RECT  6.390 3.810 6.630 4.620 ;
        RECT  5.610 4.360 6.630 4.620 ;
    END
END ad01d2

MACRO ad01d1
    CLASS CORE ;
    FOREIGN ad01d1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.823  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.630 7.470 2.870 ;
        RECT  7.230 2.090 7.470 2.870 ;
        RECT  2.860 2.630 3.300 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.648  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.120 2.020 3.860 2.390 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.036  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.980 2.100 6.870 2.390 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.300  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.170 2.580 10.520 3.650 ;
        RECT  10.170 1.550 10.410 3.650 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.071  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.660 3.330 9.220 3.570 ;
        RECT  8.970 2.220 9.220 3.570 ;
        RECT  8.460 2.220 9.220 2.460 ;
        RECT  8.460 2.020 8.960 2.460 ;
        RECT  8.720 1.420 8.960 2.460 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  9.490 4.380 9.730 5.600 ;
        RECT  8.140 4.700 8.540 5.600 ;
        RECT  4.700 4.700 5.120 5.600 ;
        RECT  3.450 4.140 3.690 5.600 ;
        RECT  0.850 4.140 1.090 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  9.460 0.000 9.700 1.420 ;
        RECT  8.010 0.000 8.250 1.280 ;
        RECT  4.870 0.000 5.110 1.280 ;
        RECT  3.450 0.000 3.690 1.340 ;
        RECT  0.820 0.000 1.060 1.240 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.170 1.630 1.880 1.870 ;
        RECT  0.150 3.600 1.910 3.840 ;
        RECT  4.040 1.620 5.820 1.860 ;
        RECT  4.390 3.130 6.060 3.370 ;
        RECT  5.820 3.130 6.060 4.120 ;
        RECT  6.100 0.980 6.500 1.840 ;
        RECT  6.100 1.600 8.110 1.840 ;
        RECT  7.870 2.800 8.700 3.040 ;
        RECT  7.870 1.600 8.110 3.420 ;
        RECT  6.360 3.180 8.110 3.420 ;
        RECT  2.250 0.980 2.490 2.350 ;
        RECT  0.120 2.110 2.490 2.350 ;
        RECT  0.120 2.110 0.360 3.360 ;
        RECT  0.120 3.120 2.480 3.360 ;
        RECT  2.240 3.660 5.580 3.900 ;
        RECT  9.690 2.390 9.930 4.050 ;
        RECT  6.390 3.810 9.930 4.050 ;
        RECT  5.340 3.660 5.580 4.600 ;
        RECT  2.240 3.120 2.480 4.540 ;
        RECT  5.340 4.360 6.630 4.600 ;
        RECT  6.390 3.810 6.630 4.620 ;
        RECT  5.610 4.360 6.630 4.620 ;
    END
END ad01d1

MACRO ad01d0
    CLASS CORE ;
    FOREIGN ad01d0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 5.600 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.823  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 2.630 7.470 2.870 ;
        RECT  7.230 2.090 7.470 2.870 ;
        RECT  2.860 2.630 3.300 3.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.648  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.120 2.080 3.860 2.390 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.036  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.980 2.100 6.870 2.390 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.696  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.170 1.650 10.520 3.890 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.696  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.660 3.570 9.220 3.810 ;
        RECT  8.970 2.230 9.220 3.810 ;
        RECT  8.460 2.020 9.070 2.460 ;
        RECT  8.670 1.620 9.070 2.460 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 4.860 10.640 5.600 ;
        RECT  9.400 4.700 9.800 5.600 ;
        RECT  8.140 4.700 8.540 5.600 ;
        RECT  4.700 4.700 5.120 5.600 ;
        RECT  3.450 4.140 3.690 5.600 ;
        RECT  0.850 4.140 1.090 5.600 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.000 10.640 0.740 ;
        RECT  9.490 0.000 9.730 1.280 ;
        RECT  8.010 0.000 8.250 1.280 ;
        RECT  4.870 0.000 5.110 1.280 ;
        RECT  3.450 0.000 3.690 1.340 ;
        RECT  0.820 0.000 1.060 1.240 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.170 1.630 1.880 1.870 ;
        RECT  0.150 3.600 1.910 3.840 ;
        RECT  4.040 1.620 5.820 1.860 ;
        RECT  4.390 3.130 6.060 3.370 ;
        RECT  5.820 3.130 6.060 4.120 ;
        RECT  6.100 0.980 6.500 1.840 ;
        RECT  6.100 1.600 8.110 1.840 ;
        RECT  7.870 2.800 8.700 3.040 ;
        RECT  7.870 1.600 8.110 3.420 ;
        RECT  6.360 3.180 8.110 3.420 ;
        RECT  2.250 0.980 2.490 2.350 ;
        RECT  0.120 2.110 2.490 2.350 ;
        RECT  0.120 2.110 0.360 3.360 ;
        RECT  0.120 3.120 2.480 3.360 ;
        RECT  2.240 3.660 5.580 3.900 ;
        RECT  5.340 3.660 5.580 4.600 ;
        RECT  6.390 4.220 9.930 4.460 ;
        RECT  9.690 2.630 9.930 4.460 ;
        RECT  2.240 3.120 2.480 4.540 ;
        RECT  5.340 4.360 6.630 4.600 ;
        RECT  5.610 4.360 6.630 4.620 ;
    END
END ad01d0

END LIBRARY

version https://git-lfs.github.com/spec/v1
oid sha256:a55187add17503f3004c7a1ce45c846afc4adc88f986cc88586e4a0be3ea0bf0
size 1736377
